----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- Description: Con RowAddr y ColAddr (que son los exponentes), se busca en la 
-- tabla de galois para la suma ---------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;

entity GaloisField_Add_5 is
generic( Bits5    : integer:=5;
         AddrBits : integer:=5);
Port
(
    Clk      : in std_logic;
    En       : in std_logic;
    RowAddr  : in std_logic_vector(AddrBits-1 downto 0);
    ColAddr  : in std_logic_vector(addrBits-1 downto 0);
    Dout     : out std_logic_vector(Bits5-1 downto 0)
);
end GaloisField_Add_5;

architecture Behavioral of GaloisField_Add_5 is
type Row is array (0 to 2**AddrBits-1) of std_logic_vector(Dout'LENGTH-1 downto 0);
type RowCol is array (0 to 2**AddrBits-1) of Row;

signal matrix : RowCol:=
(
    ("00001", "00010", "00100",	"01000", "10000", "00101",	"01010", "10100",   "01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001"),
    ("00010", "00100", "01000",	"10000", "00101", "01010",	"10100", "01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010"),
    ("00100", "01000", "10000",	"00101", "01010", "10100",	"01101", "11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100"),
    ("01000", "10000", "00101",	"01010", "10100", "01101",	"11010", "10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000"),
    ("10000", "00101", "01010",	"10100", "01101", "11010",	"10001", "00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000"),
    ("00101", "01010", "10100",	"01101", "11010", "10001",	"00111", "01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101"),
    ("01010", "10100", "01101",	"11010", "10001", "00111",	"01110", "11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010"),
    ("10100", "01101", "11010",	"10001", "00111", "01110",	"11100", "11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100"),
    ("01101", "11010", "10001",	"00111", "01110", "11100",	"11101", "11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101"),
    ("11010", "10001", "00111",	"01110", "11100", "11101",	"11111", "11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010"),
    ("10001", "00111", "01110",	"11100", "11101", "11111",	"11011", "10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001"),
    ("00111", "01110", "11100",	"11101", "11111", "11011",	"10011", "00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111"),
    ("01110", "11100", "11101",	"11111", "11011", "10011",	"00011", "00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110"),
    ("11100", "11101", "11111",	"11011", "10011", "00011",	"00110", "01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100"),
    ("11101", "11111", "11011",	"10011", "00011", "00110",	"01100", "11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101"),
    ("11111", "11011", "10011",	"00011", "00110", "01100",	"11000", "10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111"),
    ("11011", "10011", "00011",	"00110", "01100", "11000",	"10101", "01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011"),
    ("10011", "00011", "00110",	"01100", "11000", "10101",	"01111", "11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011"),
    ("00011", "00110", "01100",	"11000", "10101", "01111",	"11110", "11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011"),
    ("00110", "01100", "11000",	"10101", "01111", "11110",	"11001", "10111",	"01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110"),
    ("01100", "11000", "10101",	"01111", "11110", "11001",	"10111", "01011",	"10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100"),
    ("11000", "10101", "01111",	"11110", "11001", "10111",	"01011", "10110",	"01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000"),
    ("10101", "01111", "11110",	"11001", "10111", "01011",	"10110", "01001",	"10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101"),
    ("01111", "11110", "11001",	"10111", "01011", "10110",	"01001", "10010",	"00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111"),
    ("11110", "11001", "10111",	"01011", "10110", "01001",	"10010", "00001",	"00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110"),
    ("11001", "10111", "01011",	"10110", "01001", "10010",	"00001", "00010",	"00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001"),
    ("10111", "01011", "10110",	"01001", "10010", "00001",	"00010", "00100",	"01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111"),
    ("01011", "10110", "01001",	"10010", "00001", "00010",	"00100", "01000",	"10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011"),
    ("10110", "01001", "10010",	"00001", "00010", "00100",	"01000", "10000",	"00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110"),
    ("01001", "10010", "00001",	"00010", "00100", "01000",	"10000", "00101",	"01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001"),
    ("10010", "00001", "00010",	"00100", "01000", "10000",	"00101", "01010",	"10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010"),
    ("00001", "00010", "00100",	"01000", "10000", "00101",	"01010", "10100",	"01101",	"11010",	"10001",	"00111",	"01110",	"11100",	"11101",	"11111",	"11011",	"10011",	"00011",	"00110",	"01100",	"11000",	"10101",	"01111",	"11110",	"11001",	"10111",	"01011",	"10110",	"01001",	"10010",	"00001")
                                                                                                                                 
);
begin
process(Clk)is
begin
    if rising_edge(Clk) then
        if En ='1' then
            Dout <= matrix(conv_integer(RowAddr))(conv_integer(ColAddr));
        end if;
    end if;
end process;
--Dout <= matrix(conv_integer(RowAddr))(conv_integer(ColAddr));
end Behavioral;

library ieee;
use ieee.std_logic_1164.all;

package rom_ddm_1 is
    subtype rom_word is  std_logic_vector(5 downto 0);
    type rom_type is array (0 to 4094) of rom_word;
    constant rom_ddm1 : rom_type := (
--0
        "000001",--0
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",--10
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",--20
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",--30
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",--40
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",--50
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",--60
        "110001",
        "100001",
        "000000",
--1
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "000000",
--2
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "000000",
--3
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "000000",
--4
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "000000",
--5
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "000000",
--6
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "000000",
--7
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "000000",
--8
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "000000",
--9
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "000000",
--10
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "000000",
--11
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "000000",
--12
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "000000",
--13
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "000000",
--14
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "000000",
--15
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "000000",
--16
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "000000",
--17
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "000000",
--18
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "000000",
--19
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "000000",
--20
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "000000",
--21
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "000000",
--22
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "000000",
--23
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "000000",
--24
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "000000",
--25
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "000000",
--26
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "000000",
--27
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "000000",
--28
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "000000",
--29
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "000000",
--30
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "000000",
--31
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "000000",
--32
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "000000",
--33
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "000000",
--34
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "000000",
--35
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "000000",
--36
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "000000",
--37
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000000",
--38
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "000000",
--39
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "000000",
--40
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "000000",
--41
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "000000",
--42
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "000000",
--43
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "000000",
--44
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "000000",
--45
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "000000",
--46
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "000000",
--47
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "000000",
--48
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "000000",
--49
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "000000",
--50
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "000000",
--51
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000000",
--52
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "000000",
--53
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "000000",
--54
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "000000",
--55
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "000000",
--56
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000000",
--57
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000000",
--58
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "010000",
        "000000",
--59
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "001000",
        "000000",
--60
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000100",
        "000000",
--61
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000010",
        "000000",
--62
        "000010",
        "000100",
        "001000",
        "010000",
        "100000",
        "000011",
        "000110",
        "001100",
        "011000",
        "110000",
        "100011",
        "000101",
        "001010",
        "010100",
        "101000",
        "010011",
        "100110",
        "001111",
        "011110",
        "111100",
        "111011",
        "110101",
        "101001",
        "010001",
        "100010",
        "000111",
        "001110",
        "011100",
        "111000",
        "110011",
        "100101",
        "001001",
        "010010",
        "100100",
        "001011",
        "010110",
        "101100",
        "011011",
        "110110",
        "101111",
        "011101",
        "111010",
        "110111",
        "101101",
        "011001",
        "110010",
        "100111",
        "001101",
        "011010",
        "110100",
        "101011",
        "010101",
        "101010",
        "010111",
        "101110",
        "011111",
        "111110",
        "111111",
        "111101",
        "111001",
        "110001",
        "100001",
        "000001",
        "000000",
        others => "000000");
end rom_ddm_1;
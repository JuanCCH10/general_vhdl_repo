----------------------------------------------------------------------------------
-- Company: SEMAR
-- Engineer: TTE.FRAG.SIA.ELCO. GUILLERMO VICENCIO GUTIERREZ
-- 
-- Create Date:    12:27:30 01/03/2012 
-- Design Name:   MEMORIA
-- Module Name:    RAM_PRF - Behavioral 
-- Project Name: 
-- Target Devices: XC4VSX35-10FF668
-- Tool versions: ISE 13.1
-- Description: ALMACENAR EN EL FPGA LOS DATOS CORRESPONDIENTES A LOS NIVELES
-- DE UNA SE�AL DE FERFIL DE RANGO, ESTA SE�AL FUE MUESTREADA CON EL OSCILOSCOPIO
-- DE UN RADAR BME
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ROM_Mult_alfa is
    generic(Addrbits		: integer := 10;
			DataBits		: integer := 5
				);
	 Port (	Clk : in  STD_LOGIC;
			Addr: in  STD_LOGIC_VECTOR (Addrbits-1 downto 0);
			Rd	: in  STD_LOGIC;
			Data: out  STD_LOGIC_VECTOR (DataBits-1 downto 0));
end ROM_Mult_alfa;

architecture Behavioral of ROM_Mult_alfa is

--ROM PARA GUARDAR LOS comandos para el display oled
TYPE ROM_TYPE IS ARRAY (0 TO 2**Addrbits - 1) OF STD_LOGIC_VECTOR(DATA'range);
SIGNAL ROM: ROM_TYPE := (
33=>"00001",
34=>"00010",
36=>"00100",
40=>"01000",
48=>"10000",
37=>"00101",
42=>"01010",
52=>"10100",
45=>"01101",
58=>"11010",
49=>"10001",
39=>"00111",
46=>"01110",
60=>"11100",
61=>"11101",
63=>"11111",
59=>"11011",
51=>"10011",
35=>"00011",
38=>"00110",
44=>"01100",
56=>"11000",
53=>"10101",
47=>"01111",
62=>"11110",
57=>"11001",
55=>"10111",
43=>"01011",
54=>"10110",
41=>"01001",
50=>"10010",
--33=>"00001",
65=>"00010",
66=>"00100",
68=>"01000",
72=>"10000",
80=>"00101",
69=>"01010",
74=>"10100",
84=>"01101",
77=>"11010",
90=>"10001",
81=>"00111",
71=>"01110",
78=>"11100",
92=>"11101",
93=>"11111",
95=>"11011",
91=>"10011",
83=>"00011",
67=>"00110",
70=>"01100",
76=>"11000",
88=>"10101",
85=>"01111",
79=>"11110",
94=>"11001",
89=>"10111",
87=>"01011",
75=>"10110",
86=>"01001",
73=>"10010",
82=>"00001",
--65=>"00010",
129=>"00100",
130=>"01000",
132=>"10000",
136=>"00101",
144=>"01010",
133=>"10100",
138=>"01101",
148=>"11010",
141=>"10001",
154=>"00111",
145=>"01110",
135=>"11100",
142=>"11101",
156=>"11111",
157=>"11011",
159=>"10011",
155=>"00011",
147=>"00110",
131=>"01100",
134=>"11000",
140=>"10101",
152=>"01111",
149=>"11110",
143=>"11001",
158=>"10111",
153=>"01011",
151=>"10110",
139=>"01001",
150=>"10010",
137=>"00001",
146=>"00010",
--129=>"00100",
257=>"01000",
258=>"10000",
260=>"00101",
264=>"01010",
272=>"10100",
261=>"01101",
266=>"11010",
276=>"10001",
269=>"00111",
282=>"01110",
273=>"11100",
263=>"11101",
270=>"11111",
284=>"11011",
285=>"10011",
287=>"00011",
283=>"00110",
275=>"01100",
259=>"11000",
262=>"10101",
268=>"01111",
280=>"11110",
277=>"11001",
271=>"10111",
286=>"01011",
281=>"10110",
279=>"01001",
267=>"10010",
278=>"00001",
265=>"00010",
274=>"00100",
--257=>"01000",
513=>"10000",
514=>"00101",
516=>"01010",
520=>"10100",
528=>"01101",
517=>"11010",
522=>"10001",
532=>"00111",
525=>"01110",
538=>"11100",
529=>"11101",
519=>"11111",
526=>"11011",
540=>"10011",
541=>"00011",
543=>"00110",
539=>"01100",
531=>"11000",
515=>"10101",
518=>"01111",
524=>"11110",
536=>"11001",
533=>"10111",
527=>"01011",
542=>"10110",
537=>"01001",
535=>"10010",
523=>"00001",
534=>"00010",
521=>"00100",
530=>"01000",
--513=>"10000",
161=>"00101",
162=>"01010",
164=>"10100",
168=>"01101",
176=>"11010",
165=>"10001",
170=>"00111",
180=>"01110",
173=>"11100",
186=>"11101",
177=>"11111",
167=>"11011",
174=>"10011",
188=>"00011",
189=>"00110",
191=>"01100",
187=>"11000",
179=>"10101",
163=>"01111",
166=>"11110",
172=>"11001",
184=>"10111",
181=>"01011",
175=>"10110",
190=>"01001",
185=>"10010",
183=>"00001",
171=>"00010",
182=>"00100",
169=>"01000",
178=>"10000",
--161=>"00101",
321=>"01010",
322=>"10100",
324=>"01101",
328=>"11010",
336=>"10001",
325=>"00111",
330=>"01110",
340=>"11100",
333=>"11101",
346=>"11111",
337=>"11011",
327=>"10011",
334=>"00011",
348=>"00110",
349=>"01100",
351=>"11000",
347=>"10101",
339=>"01111",
323=>"11110",
326=>"11001",
332=>"10111",
344=>"01011",
341=>"10110",
335=>"01001",
350=>"10010",
345=>"00001",
343=>"00010",
331=>"00100",
342=>"01000",
329=>"10000",
338=>"00101",
--321=>"01010",
641=>"10100",
642=>"01101",
644=>"11010",
648=>"10001",
656=>"00111",
645=>"01110",
650=>"11100",
660=>"11101",
653=>"11111",
666=>"11011",
657=>"10011",
647=>"00011",
654=>"00110",
668=>"01100",
669=>"11000",
671=>"10101",
667=>"01111",
659=>"11110",
643=>"11001",
646=>"10111",
652=>"01011",
664=>"10110",
661=>"01001",
655=>"10010",
670=>"00001",
665=>"00010",
663=>"00100",
651=>"01000",
662=>"10000",
649=>"00101",
658=>"01010",
--641=>"10100",
417=>"01101",
418=>"11010",
420=>"10001",
424=>"00111",
432=>"01110",
421=>"11100",
426=>"11101",
436=>"11111",
429=>"11011",
442=>"10011",
433=>"00011",
423=>"00110",
430=>"01100",
444=>"11000",
445=>"10101",
447=>"01111",
443=>"11110",
435=>"11001",
419=>"10111",
422=>"01011",
428=>"10110",
440=>"01001",
437=>"10010",
431=>"00001",
446=>"00010",
441=>"00100",
439=>"01000",
427=>"10000",
438=>"00101",
425=>"01010",
434=>"10100",
--417=>"01101",
833=>"11010",
834=>"10001",
836=>"00111",
840=>"01110",
848=>"11100",
837=>"11101",
842=>"11111",
852=>"11011",
845=>"10011",
858=>"00011",
849=>"00110",
839=>"01100",
846=>"11000",
860=>"10101",
861=>"01111",
863=>"11110",
859=>"11001",
851=>"10111",
835=>"01011",
838=>"10110",
844=>"01001",
856=>"10010",
853=>"00001",
847=>"00010",
862=>"00100",
857=>"01000",
855=>"10000",
843=>"00101",
854=>"01010",
841=>"10100",
850=>"01101",
--833=>"11010",
545=>"10001",
546=>"00111",
548=>"01110",
552=>"11100",
560=>"11101",
549=>"11111",
554=>"11011",
564=>"10011",
557=>"00011",
570=>"00110",
561=>"01100",
551=>"11000",
558=>"10101",
572=>"01111",
573=>"11110",
575=>"11001",
571=>"10111",
563=>"01011",
547=>"10110",
550=>"01001",
556=>"10010",
568=>"00001",
565=>"00010",
559=>"00100",
574=>"01000",
569=>"10000",
567=>"00101",
555=>"01010",
566=>"10100",
553=>"01101",
562=>"11010",
--545=>"10001",
225=>"00111",
226=>"01110",
228=>"11100",
232=>"11101",
240=>"11111",
229=>"11011",
234=>"10011",
244=>"00011",
237=>"00110",
250=>"01100",
241=>"11000",
231=>"10101",
238=>"01111",
252=>"11110",
253=>"11001",
255=>"10111",
251=>"01011",
243=>"10110",
227=>"01001",
230=>"10010",
236=>"00001",
248=>"00010",
245=>"00100",
239=>"01000",
254=>"10000",
249=>"00101",
247=>"01010",
235=>"10100",
246=>"01101",
233=>"11010",
242=>"10001",
--225=>"00111",
449=>"01110",
450=>"11100",
452=>"11101",
456=>"11111",
464=>"11011",
453=>"10011",
458=>"00011",
468=>"00110",
461=>"01100",
474=>"11000",
465=>"10101",
455=>"01111",
462=>"11110",
476=>"11001",
477=>"10111",
479=>"01011",
475=>"10110",
467=>"01001",
451=>"10010",
454=>"00001",
460=>"00010",
472=>"00100",
469=>"01000",
463=>"10000",
478=>"00101",
473=>"01010",
471=>"10100",
459=>"01101",
470=>"11010",
457=>"10001",
466=>"00111",
--449=>"01110",
897=>"11100",
898=>"11101",
900=>"11111",
904=>"11011",
912=>"10011",
901=>"00011",
906=>"00110",
916=>"01100",
909=>"11000",
922=>"10101",
913=>"01111",
903=>"11110",
910=>"11001",
924=>"10111",
925=>"01011",
927=>"10110",
923=>"01001",
915=>"10010",
899=>"00001",
902=>"00010",
908=>"00100",
920=>"01000",
917=>"10000",
911=>"00101",
926=>"01010",
921=>"10100",
919=>"01101",
907=>"11010",
918=>"10001",
905=>"00111",
914=>"01110",
--897=>"11100",
929=>"11101",
930=>"11111",
932=>"11011",
936=>"10011",
944=>"00011",
933=>"00110",
938=>"01100",
948=>"11000",
941=>"10101",
954=>"01111",
945=>"11110",
935=>"11001",
942=>"10111",
956=>"01011",
957=>"10110",
959=>"01001",
955=>"10010",
947=>"00001",
931=>"00010",
934=>"00100",
940=>"01000",
952=>"10000",
949=>"00101",
943=>"01010",
958=>"10100",
953=>"01101",
951=>"11010",
939=>"10001",
950=>"00111",
937=>"01110",
946=>"11100",
--929=>"11101",
993=>"11111",
994=>"11011",
996=>"10011",
1000=>"00011",
1008=>"00110",
997=>"01100",
1002=>"11000",
1012=>"10101",
1005=>"01111",
1018=>"11110",
1009=>"11001",
999=>"10111",
1006=>"01011",
1020=>"10110",
1021=>"01001",
1023=>"10010",
1019=>"00001",
1011=>"00010",
995=>"00100",
998=>"01000",
1004=>"10000",
1016=>"00101",
1013=>"01010",
1007=>"10100",
1022=>"01101",
1017=>"11010",
1015=>"10001",
1003=>"00111",
1014=>"01110",
1001=>"11100",
1010=>"11101",
--993=>"11111",
865=>"11011",
866=>"10011",
868=>"00011",
872=>"00110",
880=>"01100",
869=>"11000",
874=>"10101",
884=>"01111",
877=>"11110",
890=>"11001",
881=>"10111",
871=>"01011",
878=>"10110",
892=>"01001",
893=>"10010",
895=>"00001",
891=>"00010",
883=>"00100",
867=>"01000",
870=>"10000",
876=>"00101",
888=>"01010",
885=>"10100",
879=>"01101",
894=>"11010",
889=>"10001",
887=>"00111",
875=>"01110",
886=>"11100",
873=>"11101",
882=>"11111",
--865=>"11011",
609=>"10011",
610=>"00011",
612=>"00110",
616=>"01100",
624=>"11000",
613=>"10101",
618=>"01111",
628=>"11110",
621=>"11001",
634=>"10111",
625=>"01011",
615=>"10110",
622=>"01001",
636=>"10010",
637=>"00001",
639=>"00010",
635=>"00100",
627=>"01000",
611=>"10000",
614=>"00101",
620=>"01010",
632=>"10100",
629=>"01101",
623=>"11010",
638=>"10001",
633=>"00111",
631=>"01110",
619=>"11100",
630=>"11101",
617=>"11111",
626=>"11011",
--609=>"10011",
97=>"00011",
98=>"00110",
100=>"01100",
104=>"11000",
112=>"10101",
101=>"01111",
106=>"11110",
116=>"11001",
109=>"10111",
122=>"01011",
113=>"10110",
103=>"01001",
110=>"10010",
124=>"00001",
125=>"00010",
127=>"00100",
123=>"01000",
115=>"10000",
99=>"00101",
102=>"01010",
108=>"10100",
120=>"01101",
117=>"11010",
111=>"10001",
126=>"00111",
121=>"01110",
119=>"11100",
107=>"11101",
118=>"11111",
105=>"11011",
114=>"10011",
--97=>"00011",
193=>"00110",
194=>"01100",
196=>"11000",
200=>"10101",
208=>"01111",
197=>"11110",
202=>"11001",
212=>"10111",
205=>"01011",
218=>"10110",
209=>"01001",
199=>"10010",
206=>"00001",
220=>"00010",
221=>"00100",
223=>"01000",
219=>"10000",
211=>"00101",
195=>"01010",
198=>"10100",
204=>"01101",
216=>"11010",
213=>"10001",
207=>"00111",
222=>"01110",
217=>"11100",
215=>"11101",
203=>"11111",
214=>"11011",
201=>"10011",
210=>"00011",
--193=>"00110",
385=>"01100",
386=>"11000",
388=>"10101",
392=>"01111",
400=>"11110",
389=>"11001",
394=>"10111",
404=>"01011",
397=>"10110",
410=>"01001",
401=>"10010",
391=>"00001",
398=>"00010",
412=>"00100",
413=>"01000",
415=>"10000",
411=>"00101",
403=>"01010",
387=>"10100",
390=>"01101",
396=>"11010",
408=>"10001",
405=>"00111",
399=>"01110",
414=>"11100",
409=>"11101",
407=>"11111",
395=>"11011",
406=>"10011",
393=>"00011",
402=>"00110",
--385=>"01100",
769=>"11000",
770=>"10101",
772=>"01111",
776=>"11110",
784=>"11001",
773=>"10111",
778=>"01011",
788=>"10110",
781=>"01001",
794=>"10010",
785=>"00001",
775=>"00010",
782=>"00100",
796=>"01000",
797=>"10000",
799=>"00101",
795=>"01010",
787=>"10100",
771=>"01101",
774=>"11010",
780=>"10001",
792=>"00111",
789=>"01110",
783=>"11100",
798=>"11101",
793=>"11111",
791=>"11011",
779=>"10011",
790=>"00011",
777=>"00110",
786=>"01100",
--769=>"11000",
673=>"10101",
674=>"01111",
676=>"11110",
680=>"11001",
688=>"10111",
677=>"01011",
682=>"10110",
692=>"01001",
685=>"10010",
698=>"00001",
689=>"00010",
679=>"00100",
686=>"01000",
700=>"10000",
701=>"00101",
703=>"01010",
699=>"10100",
691=>"01101",
675=>"11010",
678=>"10001",
684=>"00111",
696=>"01110",
693=>"11100",
687=>"11101",
702=>"11111",
697=>"11011",
695=>"10011",
683=>"00011",
694=>"00110",
681=>"01100",
690=>"11000",
--673=>"10101",
481=>"01111",
482=>"11110",
484=>"11001",
488=>"10111",
496=>"01011",
485=>"10110",
490=>"01001",
500=>"10010",
493=>"00001",
506=>"00010",
497=>"00100",
487=>"01000",
494=>"10000",
508=>"00101",
509=>"01010",
511=>"10100",
507=>"01101",
499=>"11010",
483=>"10001",
486=>"00111",
492=>"01110",
504=>"11100",
501=>"11101",
495=>"11111",
510=>"11011",
505=>"10011",
503=>"00011",
491=>"00110",
502=>"01100",
489=>"11000",
498=>"10101",
--481=>"01111",
961=>"11110",
962=>"11001",
964=>"10111",
968=>"01011",
976=>"10110",
965=>"01001",
970=>"10010",
980=>"00001",
973=>"00010",
986=>"00100",
977=>"01000",
967=>"10000",
974=>"00101",
988=>"01010",
989=>"10100",
991=>"01101",
987=>"11010",
979=>"10001",
963=>"00111",
966=>"01110",
972=>"11100",
984=>"11101",
981=>"11111",
975=>"11011",
990=>"10011",
985=>"00011",
983=>"00110",
971=>"01100",
982=>"11000",
969=>"10101",
978=>"01111",
--961=>"11110",
801=>"11001",
802=>"10111",
804=>"01011",
808=>"10110",
816=>"01001",
805=>"10010",
810=>"00001",
820=>"00010",
813=>"00100",
826=>"01000",
817=>"10000",
807=>"00101",
814=>"01010",
828=>"10100",
829=>"01101",
831=>"11010",
827=>"10001",
819=>"00111",
803=>"01110",
806=>"11100",
812=>"11101",
824=>"11111",
821=>"11011",
815=>"10011",
830=>"00011",
825=>"00110",
823=>"01100",
811=>"11000",
822=>"10101",
809=>"01111",
818=>"11110",
--801=>"11001",
737=>"10111",
738=>"01011",
740=>"10110",
744=>"01001",
752=>"10010",
741=>"00001",
746=>"00010",
756=>"00100",
749=>"01000",
762=>"10000",
753=>"00101",
743=>"01010",
750=>"10100",
764=>"01101",
765=>"11010",
767=>"10001",
763=>"00111",
755=>"01110",
739=>"11100",
742=>"11101",
748=>"11111",
760=>"11011",
757=>"10011",
751=>"00011",
766=>"00110",
761=>"01100",
759=>"11000",
747=>"10101",
758=>"01111",
745=>"11110",
754=>"11001",
--737=>"10111",
353=>"01011",
354=>"10110",
356=>"01001",
360=>"10010",
368=>"00001",
357=>"00010",
362=>"00100",
372=>"01000",
365=>"10000",
378=>"00101",
369=>"01010",
359=>"10100",
366=>"01101",
380=>"11010",
381=>"10001",
383=>"00111",
379=>"01110",
371=>"11100",
355=>"11101",
358=>"11111",
364=>"11011",
376=>"10011",
373=>"00011",
367=>"00110",
382=>"01100",
377=>"11000",
375=>"10101",
363=>"01111",
374=>"11110",
361=>"11001",
370=>"10111",
--353=>"01011",
705=>"10110",
706=>"01001",
708=>"10010",
712=>"00001",
720=>"00010",
709=>"00100",
714=>"01000",
724=>"10000",
717=>"00101",
730=>"01010",
721=>"10100",
711=>"01101",
718=>"11010",
732=>"10001",
733=>"00111",
735=>"01110",
731=>"11100",
723=>"11101",
707=>"11111",
710=>"11011",
716=>"10011",
728=>"00011",
725=>"00110",
719=>"01100",
734=>"11000",
729=>"10101",
727=>"01111",
715=>"11110",
726=>"11001",
713=>"10111",
722=>"01011",
--705=>"10110",
289=>"01001",
290=>"10010",
292=>"00001",
296=>"00010",
304=>"00100",
293=>"01000",
298=>"10000",
308=>"00101",
301=>"01010",
314=>"10100",
305=>"01101",
295=>"11010",
302=>"10001",
316=>"00111",
317=>"01110",
319=>"11100",
315=>"11101",
307=>"11111",
291=>"11011",
294=>"10011",
300=>"00011",
312=>"00110",
309=>"01100",
303=>"11000",
318=>"10101",
313=>"01111",
311=>"11110",
299=>"11001",
310=>"10111",
297=>"01011",
306=>"10110",
--289=>"01001",
577=>"10010",
578=>"00001",
580=>"00010",
584=>"00100",
592=>"01000",
581=>"10000",
586=>"00101",
596=>"01010",
589=>"10100",
602=>"01101",
593=>"11010",
583=>"10001",
590=>"00111",
604=>"01110",
605=>"11100",
607=>"11101",
603=>"11111",
595=>"11011",
579=>"10011",
582=>"00011",
588=>"00110",
600=>"01100",
597=>"11000",
591=>"10101",
606=>"01111",
601=>"11110",
599=>"11001",
587=>"10111",
598=>"01011",
585=>"10110",
594=>"01001",
--577=>"10010",
--33=>"00001",
--34=>"00010",
--36=>"00100",
--40=>"01000",
--48=>"10000",
--37=>"00101",
--42=>"01010",
--52=>"10100",
--45=>"01101",
--58=>"11010",
--49=>"10001",
--39=>"00111",
--46=>"01110",
--60=>"11100",
--61=>"11101",
--63=>"11111",
--59=>"11011",
--51=>"10011",
--35=>"00011",
--38=>"00110",
--44=>"01100",
--56=>"11000",
--53=>"10101",
--47=>"01111",
--62=>"11110",
--57=>"11001",
--55=>"10111",
--43=>"01011",
--54=>"10110",
--41=>"01001",
--50=>"10010",
--33=>"00001",

others=>"00000");
begin

process(clk)  begin
	if rising_edge(clk)  then
		if Rd = '1' then
			Data <= rom(conv_integer(addr));  -- First register
		end if;
	end if;
end process;
end Behavioral;


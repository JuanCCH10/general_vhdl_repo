library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity prod_alpha_tb is
end prod_alpha_tb;

architecture Behavioral of prod_alpha_tb is

    component prod_alpha is
        Port (
            alphaA : in std_logic_vector(5 downto 0);
            alphaB : in std_logic_vector(5 downto 0);
            alphaR : out std_logic_vector(5 downto 0)
        );
    end component;
    
    constant per : time := 10ns;
    signal clk : std_logic;
    signal alphaA, alphaB, alphaR : std_logic_vector(5 downto 0);

begin

    clk_gen : process is begin
        clk <= '1';
        wait for per/2;
        clk <= '0';
        wait for per/2;
    end process;
    
    conexiones : prod_alpha
    port map(
        alphaA => alphaA,
        alphaB => alphaB,
        alphaR => alphaR
    );
    
    estimulos : process is begin
        alphaA <= "000000";
        alphaB <= "000000";
        wait for per;
        alphaA <= "000000";
        alphaB <= "000001";
        wait for per;
        alphaA <= "000001";
        alphaB <= "000000";
        wait for per;
        alphaA <= "000001";
        alphaB <= "000001";
        wait for per;
        alphaA <= "000010";
        alphaB <= "000001";
        wait for per;
        alphaA <= "000100";
        alphaB <= "000001";
        wait for per;
        alphaA <= "001000";
        alphaB <= "000001";
        wait for per;
        alphaA <= "010000";
        alphaB <= "000001";
        wait for per;
        alphaA <= "100000";
        alphaB <= "000001";
        wait for per;
        alphaA <= "000011";
        alphaB <= "000001";
        wait for per;
        alphaA <= "000110";
        alphaB <= "000001";
        wait for per;
        alphaA <= "001100";
        alphaB <= "000001";
        wait for per;
        alphaA <= "011000";
        alphaB <= "000001";
        wait for per;
        alphaA <= "110000";
        alphaB <= "000001";
        wait for per;
        alphaA <= "100011";
        alphaB <= "000001";
        wait for per;
        alphaA <= "000101";
        alphaB <= "000001";
        wait for per;
        alphaA <= "001010";
        alphaB <= "000001";
        wait for per;
        alphaA <= "010100";
        alphaB <= "000001";
        wait for per;
        alphaA <= "101000";
        alphaB <= "000001";
        wait for per;
        alphaA <= "010011";
        alphaB <= "000001";
        wait for per;
        alphaA <= "100110";
        alphaB <= "000001";
        wait for per;
        alphaA <= "001111";
        alphaB <= "000001";
        wait for per;
        alphaA <= "011110";
        alphaB <= "000001";
        wait for per;
        alphaA <= "111100";
        alphaB <= "000001";
        wait for per;
        alphaA <= "111011";
        alphaB <= "000001";
        wait for per;
        alphaA <= "110101";
        alphaB <= "000001";
        wait for per;
        alphaA <= "101001";
        alphaB <= "000001";
        wait for per;
        alphaA <= "010001";
        alphaB <= "000001";
        wait for per;
        alphaA <= "100010";
        alphaB <= "000001";
        wait for per;
        alphaA <= "000111";
        alphaB <= "000001";
        wait for per;
        alphaA <= "001110";
        alphaB <= "000001";
        wait for per;
        alphaA <= "011100";
        alphaB <= "000001";
        wait for per;
        alphaA <= "111000";
        alphaB <= "000001";
        wait for per;
        alphaA <= "110011";
        alphaB <= "000001";
        wait for per;
        alphaA <= "100101";
        alphaB <= "000001";
        wait for per;
        alphaA <= "001001";
        alphaB <= "000001";
        wait for per;
        alphaA <= "010010";
        alphaB <= "000001";
        wait for per;
        alphaA <= "100100";
        alphaB <= "000001";
        wait for per;
        alphaA <= "001011";
        alphaB <= "000001";
        wait for per;
        alphaA <= "010110";
        alphaB <= "000001";
        wait for per;
        alphaA <= "101100";
        alphaB <= "000001";
        wait for per;
        alphaA <= "011011";
        alphaB <= "000001";
        wait for per;
        alphaA <= "110110";
        alphaB <= "000001";
        wait for per;
        alphaA <= "101111";
        alphaB <= "000001";
        wait for per;
        alphaA <= "011101";
        alphaB <= "000001";
        wait for per;
        alphaA <= "111010";
        alphaB <= "000001";
        wait for per;
        alphaA <= "110111";
        alphaB <= "000001";
        wait for per;
        alphaA <= "101101";
        alphaB <= "000001";
        wait for per;
        alphaA <= "011001";
        alphaB <= "000001";
        wait for per;
        alphaA <= "110010";
        alphaB <= "000001";
        wait for per;
        alphaA <= "100111";
        alphaB <= "000001";
        wait for per;
        alphaA <= "001101";
        alphaB <= "000001";
        wait for per;
        alphaA <= "011010";
        alphaB <= "000001";
        wait for per;
        alphaA <= "110100";
        alphaB <= "000001";
        wait for per;
        alphaA <= "101011";
        alphaB <= "000001";
        wait for per;
        alphaA <= "010101";
        alphaB <= "000001";
        wait for per;
        alphaA <= "101010";
        alphaB <= "000001";
        wait for per;
        alphaA <= "010111";
        alphaB <= "000001";
        wait for per;
        alphaA <= "101110";
        alphaB <= "000001";
        wait for per;
        alphaA <= "011111";
        alphaB <= "000001";
        wait for per;
        alphaA <= "111110";
        alphaB <= "000001";
        wait for per;
        alphaA <= "111111";
        alphaB <= "000001";
        wait for per;
        alphaA <= "111101";
        alphaB <= "000001";
        wait for per;
        alphaA <= "111001";
        alphaB <= "000001";
        wait for per;
        alphaA <= "110001";
        alphaB <= "000001";
        wait for per;
        alphaA <= "100001";
        alphaB <= "000001";
        wait for 3*per;


        alphaA <= "000000";
        alphaB <= "000010";
        wait for per;
        alphaA <= "000001";
        alphaB <= "000010";
        wait for per;
        alphaA <= "000010";
        alphaB <= "000010";
        wait for per;
        alphaA <= "000100";
        alphaB <= "000010";
        wait for per;
        alphaA <= "001000";
        alphaB <= "000010";
        wait for per;
        alphaA <= "010000";
        alphaB <= "000010";
        wait for per;
        alphaA <= "100000";
        alphaB <= "000010";
        wait for per;
        alphaA <= "000011";
        alphaB <= "000010";
        wait for per;
        alphaA <= "000110";
        alphaB <= "000010";
        wait for per;
        alphaA <= "001100";
        alphaB <= "000010";
        wait for per;
        alphaA <= "011000";
        alphaB <= "000010";
        wait for per;
        alphaA <= "110000";
        alphaB <= "000010";
        wait for per;
        alphaA <= "100011";
        alphaB <= "000010";
        wait for per;
        alphaA <= "000101";
        alphaB <= "000010";
        wait for per;
        alphaA <= "001010";
        alphaB <= "000010";
        wait for per;
        alphaA <= "010100";
        alphaB <= "000010";
        wait for per;
        alphaA <= "101000";
        alphaB <= "000010";
        wait for per;
        alphaA <= "010011";
        alphaB <= "000010";
        wait for per;
        alphaA <= "100110";
        alphaB <= "000010";
        wait for per;
        alphaA <= "001111";
        alphaB <= "000010";
        wait for per;
        alphaA <= "011110";
        alphaB <= "000010";
        wait for per;
        alphaA <= "111100";
        alphaB <= "000010";
        wait for per;
        alphaA <= "111011";
        alphaB <= "000010";
        wait for per;
        alphaA <= "110101";
        alphaB <= "000010";
        wait for per;
        alphaA <= "101001";
        alphaB <= "000010";
        wait for per;
        alphaA <= "010001";
        alphaB <= "000010";
        wait for per;
        alphaA <= "100010";
        alphaB <= "000010";
        wait for per;
        alphaA <= "000111";
        alphaB <= "000010";
        wait for per;
        alphaA <= "001110";
        alphaB <= "000010";
        wait for per;
        alphaA <= "011100";
        alphaB <= "000010";
        wait for per;
        alphaA <= "111000";
        alphaB <= "000010";
        wait for per;
        alphaA <= "110011";
        alphaB <= "000010";
        wait for per;
        alphaA <= "100101";
        alphaB <= "000010";
        wait for per;
        alphaA <= "001001";
        alphaB <= "000010";
        wait for per;
        alphaA <= "010010";
        alphaB <= "000010";
        wait for per;
        alphaA <= "100100";
        alphaB <= "000010";
        wait for per;
        alphaA <= "001011";
        alphaB <= "000010";
        wait for per;
        alphaA <= "010110";
        alphaB <= "000010";
        wait for per;
        alphaA <= "101100";
        alphaB <= "000010";
        wait for per;
        alphaA <= "011011";
        alphaB <= "000010";
        wait for per;
        alphaA <= "110110";
        alphaB <= "000010";
        wait for per;
        alphaA <= "101111";
        alphaB <= "000010";
        wait for per;
        alphaA <= "011101";
        alphaB <= "000010";
        wait for per;
        alphaA <= "111010";
        alphaB <= "000010";
        wait for per;
        alphaA <= "110111";
        alphaB <= "000010";
        wait for per;
        alphaA <= "101101";
        alphaB <= "000010";
        wait for per;
        alphaA <= "011001";
        alphaB <= "000010";
        wait for per;
        alphaA <= "110010";
        alphaB <= "000010";
        wait for per;
        alphaA <= "100111";
        alphaB <= "000010";
        wait for per;
        alphaA <= "001101";
        alphaB <= "000010";
        wait for per;
        alphaA <= "011010";
        alphaB <= "000010";
        wait for per;
        alphaA <= "110100";
        alphaB <= "000010";
        wait for per;
        alphaA <= "101011";
        alphaB <= "000010";
        wait for per;
        alphaA <= "010101";
        alphaB <= "000010";
        wait for per;
        alphaA <= "101010";
        alphaB <= "000010";
        wait for per;
        alphaA <= "010111";
        alphaB <= "000010";
        wait for per;
        alphaA <= "101110";
        alphaB <= "000010";
        wait for per;
        alphaA <= "011111";
        alphaB <= "000010";
        wait for per;
        alphaA <= "111110";
        alphaB <= "000010";
        wait for per;
        alphaA <= "111111";
        alphaB <= "000010";
        wait for per;
        alphaA <= "111101";
        alphaB <= "000010";
        wait for per;
        alphaA <= "111001";
        alphaB <= "000010";
        wait for per;
        alphaA <= "110001";
        alphaB <= "000010";
        wait for per;
        alphaA <= "100001";
        alphaB <= "000010";
        wait;
    end process;
end Behavioral;

----------------------------------------------------------------------------------
-- Company: SEMAR
-- Engineer: TTE.FRAG.SIA.ELCO. GUILLERMO VICENCIO GUTIERREZ
-- 
-- Create Date:    19:27:30 19/11/2021
-- Design Name:   MEMORIA
-- Module Name:    ROM_Conf_CML - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: Vivado
-- Description: 
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ROM_Simbolos_dam_r41 is
    generic(Addrbits		: integer := 6;
				DataBits		: integer := 8
				);
	 Port ( Clk : in  STD_LOGIC;
			  Addr: in  STD_LOGIC_VECTOR (Addrbits-1 downto 0);
           Rd	: in  STD_LOGIC;
			  Data: out  STD_LOGIC_VECTOR (DataBits-1 downto 0));
end ROM_Simbolos_dam_r41;

architecture Behavioral of ROM_Simbolos_dam_r41 is

--ROM PARA GUARDAR LOS comandos para el display oled
TYPE ROM_TYPE IS ARRAY (0 TO 2**Addrbits - 1) OF STD_LOGIC_VECTOR(DATA'range);
SIGNAL ROM: ROM_TYPE := (
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"00",
"00",
"00",
"00",
"11",
"00",
"11",
"00",
"11",
"10",
"11",
"01",
"01",
"11",
"01",
"11",
"11",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"00",
"11",
"01",
"11",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"11",
"10",
"10",
"11",
"01",
"01",
"11",
"10",
"00",
"00",
"10",
"01",
"01",
"00",
"01",
"01",
"00",
"10",
"01",
"11",
"11",
"00",
"00",
"10",
"10",
"10",
"00",
"10",
"00",
"11",
"01",
"01",
"01",
"00",
"00",
"00",
"11",
"01",
"10",
"01",
"11",
"11",
"00",
"11",
"01",
"00",
"01",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"11",
"01",
"01",
"00",
"00",
"01",
"11",
"10",
"01",
"00",
"00",
"10",
"00",
"01",
"11",
"10",
"10",
"10",
"00",
"10",
"00",
"11",
"01",
"01",
"10",
"00",
"10",
"11",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"01",
"00",
"10",
"10",
"10",
"01",
"01",
"11",
"10",
"00",
"11",
"01",
"11",
"00",
"01",
"10",
"00",
"01",
"00",
"10",
"10",
"10",
"01",
"01",
"10",
"01",
"01",
"00",
"01",
"10",
"11",
"10",
"00",
"00",
"11",
"00",
"00",
"10",
"10",
"01",
"00",
"11",
"11",
"10",
"00",
"00",
"00",
"11",
"00",
"01",
"11",
"01",
"01",
"01",
"00",
"11",
"00",
"01",
"11",
"01",
"01",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"10",
"01",
"11",
"11",
"00",
"00",
"10",
"00",
"01",
"10",
"10",
"01",
"01",
"00",
"00",
"00",
"00",
"11",
"10",
"10",
"00",
"10",
"00",
"01",
"01",
"10",
"00",
"11",
"10",
"00",
"00",
"00",
"10",
"00",
"01",
"01",
"11",
"01",
"00",
"11",
"01",
"10",
"01",
"10",
"11",
"00",
"00",
"01",
"11",
"10",
"00",
"01",
"01",
"11",
"00",
"10",
"01",
"11",
"01",
"10",
"01",
"11",
"00",
"00",
"10",
"11",
"01",
"01",
"10",
"10",
"00",
"00",
"11",
"01",
"10",
"01",
"11",
"01",
"01",
"11",
"00",
"01",
"11",
"01",
"00",
"00",
"00",
"00",
"01",
"11",
"10",
"00",
"11",
"01",
"01",
"10",
"00",
"11",
"00",
"00",
"10",
"11",
"00",
"10",
"11",
"11",
"00",
"11",
"01",
"10",
"00",
"10",
"11",
"11",
"11",
"11",
"10",
"00",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"00",
"11",
"00",
"01",
"01",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"01",
"00",
"11",
"10",
"00",
"10",
"11",
"00",
"01",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"00",
"00",
"11",
"01",
"11",
"10",
"00",
"10",
"00",
"10",
"01",
"01",
"11",
"01",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"00",
"01",
"01",
"11",
"11",
"11",
"00",
"11",
"00",
"10",
"01",
"11",
"11",
"01",
"00",
"00",
"00",
"11",
"10",
"11",
"01",
"00",
"01",
"10",
"11",
"10",
"11",
"00",
"01",
"10",
"00",
"11",
"00",
"11",
"11",
"01",
"01",
"11",
"10",
"10",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"01",
"00",
"00",
"11",
"10",
"01",
"11",
"11",
"10",
"10",
"11",
"11",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"00",
"11",
"10",
"00",
"01",
"00",
"11",
"10",
"01",
"11",
"11",
"10",
"01",
"00",
"00",
"11",
"11",
"11",
"01",
"11",
"01",
"10",
"01",
"01",
"10",
"11",
"01",
"00",
"00",
"01",
"11",
"01",
"10",
"00",
"11",
"10",
"10",
"01",
"11",
"01",
"11",
"11",
"10",
"01",
"10",
"01",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"00",
"00",
"11",
"11",
"11",
"10",
"11",
"10",
"10",
"11",
"01",
"01",
"00",
"10",
"00",
"00",
"11",
"01",
"01",
"11",
"10",
"11",
"00",
"10",
"00",
"11",
"00",
"00",
"10",
"01",
"11",
"10",
"11",
"10",
"00",
"01",
"11",
"00",
"11",
"01",
"01",
"00",
"11",
"00",
"10",
"11",
"01",
"01",
"01",
"11",
"01",
"00",
"11",
"11",
"11",
"11",
"11",
"00",
"01",
"00",
"01",
"10",
"11",
"00",
"01",
"10",
"11",
"10",
"10",
"11",
"11",
"10",
"11",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"00",
"11",
"00",
"10",
"11",
"01",
"11",
"11",
"10",
"01",
"11",
"01",
"00",
"01",
"10",
"00",
"11",
"01",
"00",
"11",
"11",
"10",
"10",
"01",
"01",
"10",
"00",
"00",
"00",
"11",
"01",
"10",
"10",
"11",
"00",
"01",
"01",
"10",
"10",
"11",
"11",
"11",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"01",
"11",
"00",
"11",
"00",
"01",
"11",
"00",
"10",
"10",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"00",
"10",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"01",
"10",
"01",
"01",
"11",
"11",
"00",
"10",
"00",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"01",
"10",
"01",
"00",
"10",
"00",
"10",
"10",
"01",
"10",
"10",
"10",
"10",
"11",
"00",
"00",
"10",
"01",
"11",
"00",
"00",
"10",
"10",
"11",
"10",
"00",
"11",
"00",
"00",
"10",
"11",
"11",
"00",
"01",
"00",
"11",
"10",
"00",
"01",
"01",
"11",
"01",
"00",
"00",
"10",
"00",
"10",
"00",
"01",
"00",
"10",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"10",
"11",
"10",
"10",
"11",
"10",
"11",
"00",
"00",
"00",
"10",
"11",
"00",
"00",
"01",
"00",
"01",
"10",
"11",
"11",
"00",
"11",
"01",
"10",
"01",
"10",
"11",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"10",
"00",
"10",
"11",
"01",
"10",
"00",
"10",
"01",
"10",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"10",
"01",
"01",
"10",
"10",
"00",
"10",
"11",
"11",
"10",
"01",
"00",
"00",
"11",
"00",
"10",
"00",
"00",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"00",
"00",
"00",
"10",
"00",
"01",
"00",
"00",
"01",
"00",
"11",
"00",
"11",
"11",
"10",
"01",
"01",
"10",
"10",
"01",
"00",
"00",
"10",
"10",
"00",
"11",
"10",
"01",
"11",
"11",
"11",
"00",
"00",
"01",
"00",
"11",
"10",
"10",
"10",
"10",
"10",
"11",
"01",
"11",
"00",
"10",
"11",
"10",
"11",
"01",
"00",
"01",
"00",
"10",
"00",
"11",
"11",
"10",
"10",
"00",
"11",
"00",
"00",
"01",
"11",
"11",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"10",
"00",
"00",
"01",
"11",
"11",
"10",
"10",
"11",
"01",
"00",
"01",
"10",
"00",
"00",
"00",
"11",
"11",
"10",
"11",
"11",
"11",
"11",
"00",
"10",
"00",
"01",
"00",
"10",
"00",
"00",
"11",
"11",
"00",
"00",
"00",
"11",
"10",
"01",
"11",
"00",
"01",
"00",
"10",
"01",
"10",
"00",
"01",
"11",
"00",
"01",
"10",
"01",
"01",
"10",
"00",
"01",
"11",
"00",
"11",
"11",
"01",
"10",
"11",
"11",
"11",
"00",
"01",
"10",
"01",
"00",
"11",
"01",
"10",
"11",
"00",
"01",
"11",
"10",
"00",
"01",
"00",
"01",
"10",
"00",
"00",
"01",
"01",
"11",
"10",
"01",
"01",
"00",
"10",
"11",
"11",
"01",
"01",
"10",
"11",
"00",
"10",
"01",
"00",
"01",
"10",
"11",
"11",
"01",
"01",
"10",
"01",
"11",
"10",
"00",
"01",
"11",
"00",
"10",
"01",
"10",
"00",
"00",
"11",
"11",
"11",
"00",
"01",
"10",
"11",
"00",
"11",
"11",
"10",
"00",
"00",
"10",
"01",
"00",
"01",
"11",
"00",
"00",
"11",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"01",
"01",
"00",
"00",
"00",
"01",
"11",
"10",
"00",
"11",
"00",
"01",
"10",
"01",
"00",
"00",
"11",
"00",
"11",
"11",
"01",
"01",
"11",
"01",
"10",
"00",
"10",
"00",
"01",
"01",
"00",
"10",
"00",
"01",
"00",
"01",
"00",
"00",
"10",
"01",
"10",
"11",
"10",
"10",
"10",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"10",
"00",
"11",
"00",
"11",
"01",
"01",
"10",
"11",
"00",
"10",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"00",
"01",
"00",
"11",
"00",
"00",
"00",
"11",
"11",
"01",
"00",
"11",
"10",
"00",
"00",
"11",
"10",
"00",
"11",
"01",
"11",
"01",
"10",
"10",
"01",
"10",
"01",
"11",
"01",
"01",
"10",
"11",
"11",
"10",
"10",
"11",
"00",
"10",
"01",
"01",
"01",
"01",
"10",
"10",
"01",
"11",
"11",
"01",
"01",
"10",
"11",
"11",
"00",
"11",
"11",
"01",
"11",
"11",
"00",
"11",
"01",
"10",
"01",
"11",
"10",
"01",
"10",
"11",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"01",
"01",
"11",
"11",
"01",
"10",
"10",
"11",
"01",
"11",
"01",
"00",
"10",
"11",
"00",
"10",
"00",
"01",
"10",
"01",
"01",
"01",
"10",
"10",
"00",
"01",
"00",
"11",
"10",
"11",
"01",
"10",
"01",
"01",
"10",
"10",
"11",
"11",
"11",
"10",
"01",
"11",
"11",
"10",
"01",
"01",
"01",
"00",
"10",
"00",
"00",
"00",
"11",
"10",
"01",
"00",
"11",
"11",
"01",
"01",
"00",
"00",
"00",
"11",
"00",
"11",
"11",
"11",
"00",
"00",
"01",
"11",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"01",
"11",
"00",
"01",
"01",
"10",
"01",
"01",
"00",
"10",
"01",
"01",
"01",
"10",
"10",
"10",
"11",
"01",
"11",
"11",
"10",
"11",
"01",
"00",
"10",
"01",
"10",
"00",
"11",
"00",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"00",
"00",
"01",
"10",
"11",
"01",
"11",
"00",
"01",
"10",
"10",
"11",
"11",
"11",
"10",
"10",
"01",
"11",
"11",
"10",
"10",
"00",
"01",
"00",
"10",
"11",
"00",
"00",
"11",
"10",
"11",
"10",
"11",
"01",
"01",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"10",
"01",
"00",
"01",
"11",
"00",
"00",
"01",
"10",
"11",
"00",
"01",
"00",
"10",
"11",
"10",
"11",
"01",
"10",
"11",
"11",
"01",
"01",
"00",
"00",
"11",
"10",
"10",
"10",
"10",
"00",
"11",
"10",
"01",
"00",
"11",
"01",
"00",
"11",
"11",
"00",
"11",
"00",
"11",
"11",
"01",
"10",
"01",
"11",
"11",
"01",
"11",
"10",
"00",
"00",
"01",
"00",
"01",
"00",
"01",
"11",
"00",
"11",
"01",
"10",
"11",
"11",
"00",
"10",
"10",
"01",
"01",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"00",
"01",
"11",
"01",
"11",
"11",
"10",
"00",
"01",
"11",
"11",
"01",
"00",
"10",
"10",
"10",
"10",
"01",
"10",
"00",
"00",
"11",
"10",
"00",
"10",
"01",
"11",
"00",
"01",
"10",
"00",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"10",
"01",
"01",
"00",
"10",
"10",
"10",
"00",
"01",
"11",
"00",
"00",
"10",
"10",
"00",
"00",
"01",
"11",
"00",
"11",
"00",
"00",
"00",
"10",
"01",
"11",
"10",
"10",
"01",
"01",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"10",
"10",
"01",
"01",
"10",
"11",
"10",
"10",
"01",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"01",
"10",
"00",
"11",
"10",
"11",
"10",
"00",
"11",
"10",
"10",
"11",
"11",
"01",
"11",
"11",
"11",
"00",
"10",
"01",
"10",
"10",
"10",
"11",
"10",
"11",
"10",
"01",
"11",
"01",
"10",
"01",
"10",
"10",
"11",
"01",
"10",
"10",
"11",
"00",
"11",
"11",
"00",
"00",
"00",
"10",
"01",
"01",
"01",
"11",
"01",
"01",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"00",
"10",
"00",
"10",
"10",
"00",
"00",
"00",
"11",
"10",
"10",
"10",
"11",
"11",
"10",
"01",
"01",
"11",
"11",
"00",
"01",
"10",
"00",
"10",
"10",
"01",
"11",
"11",
"10",
"11",
"01",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"11",
"11",
"01",
"10",
"00",
"00",
"11",
"11",
"00",
"10",
"00",
"11",
"10",
"10",
"00",
"01",
"10",
"11",
"10",
"11",
"00",
"10",
"00",
"10",
"01",
"01",
"11",
"11",
"10",
"10",
"11",
"10",
"11",
"10",
"11",
"11",
"00",
"00",
"01",
"01",
"00",
"00",
"11",
"10",
"10",
"00",
"01",
"10",
"10",
"11",
"01",
"01",
"11",
"01",
"01",
"10",
"10",
"00",
"00",
"10",
"10",
"11",
"01",
"10",
"11",
"00",
"10",
"01",
"11",
"11",
"01",
"11",
"01",
"10",
"01",
"11",
"00",
"01",
"00",
"10",
"10",
"11",
"10",
"01",
"11",
"11",
"00",
"00",
"11",
"01",
"01",
"11",
"10",
"10",
"01",
"10",
"10",
"01",
"11",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"00",
"00",
"11",
"10",
"10",
"01",
"00",
"00",
"10",
"01",
"01",
"11",
"01",
"10",
"00",
"11",
"11",
"11",
"01",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"00",
"01",
"00",
"10",
"10",
"00",
"00",
"10",
"10",
"00",
"11",
"11",
"00",
"11",
"01",
"00",
"00",
"00",
"01",
"10",
"00",
"00",
"10",
"11",
"10",
"11",
"11",
"11",
"11",
"10",
"10",
"11",
"01",
"10",
"00",
"01",
"00",
"00",
"00",
"00",
"10",
"01",
"10",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"00",
"10",
"00",
"00",
"10",
"10",
"11",
"01",
"01",
"01",
"11",
"10",
"11",
"10",
"10",
"10",
"01",
"00",
"00",
"00",
"10",
"01",
"00",
"10",
"10",
"01",
"00",
"10",
"01",
"01",
"11",
"01",
"10",
"11",
"00",
"10",
"10",
"01",
"00",
"01",
"10",
"10",
"00",
"01",
"01",
"01",
"10",
"11",
"10",
"01",
"00",
"10",
"10",
"01",
"10",
"00",
"01",
"01",
"10",
"01",
"01",
"00",
"00",
"10",
"01",
"00",
"10",
"11",
"01",
"01",
"00",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"00",
"00",
"10",
"00",
"00",
"00",
"11",
"01",
"00",
"10",
"01",
"10",
"11",
"00",
"00",
"10",
"01",
"01",
"11",
"01",
"01",
"10",
"01",
"10",
"01",
"11",
"01",
"11",
"01",
"10",
"10",
"10",
"00",
"10",
"01",
"00",
"00",
"00",
"11",
"01",
"10",
"10",
"01",
"10",
"00",
"11",
"01",
"11",
"00",
"00",
"00",
"01",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"11",
"11",
"00",
"00",
"00",
"11",
"11",
"00",
"00",
"10",
"01",
"11",
"10",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"11",
"10",
"01",
"11",
"00",
"00",
"00",
"10",
"01",
"10",
"11",
"00",
"01",
"00",
"00",
"10",
"11",
"11",
"10",
"11",
"01",
"00",
"10",
"10",
"01",
"01",
"00",
"11",
"00",
"11",
"10",
"11",
"11",
"01",
"01",
"01",
"00",
"00",
"11",
"01",
"00",
"01",
"01",
"10",
"10",
"10",
"00",
"01",
"00",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"10",
"10",
"11",
"11",
"01",
"01",
"01",
"00",
"00",
"01",
"10",
"11",
"10",
"00",
"00",
"00",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"10",
"00",
"00",
"01",
"11",
"01",
"00",
"00",
"11",
"10",
"01",
"01",
"00",
"00",
"11",
"01",
"10",
"10",
"11",
"10",
"11",
"11",
"11",
"11",
"01",
"11",
"00",
"11",
"10",
"11",
"10",
"00",
"01",
"00",
"01",
"01",
"11",
"11",
"10",
"00",
"01",
"01",
"11",
"00",
"01",
"01",
"01",
"11",
"01",
"10",
"01",
"00",
"01",
"11",
"10",
"10",
"10",
"10",
"01",
"11",
"00",
"00",
"10",
"11",
"00",
"11",
"00",
"10",
"01",
"11",
"01",
"10",
"10",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"11",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"00",
"01",
"00",
"10",
"10",
"10",
"11",
"10",
"00",
"11",
"01",
"11",
"10",
"10",
"10",
"00",
"00",
"10",
"10",
"01",
"00",
"10",
"10",
"01",
"11",
"01",
"10",
"11",
"01",
"11",
"10",
"01",
"01",
"01",
"01",
"01",
"10",
"11",
"11",
"00",
"10",
"01",
"11",
"01",
"00",
"11",
"11",
"11",
"10",
"01",
"00",
"01",
"10",
"01",
"00",
"11",
"10",
"00",
"00",
"11",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"11",
"01",
"00",
"01",
"11",
"10",
"11",
"01",
"11",
"00",
"00",
"10",
"10",
"00",
"11",
"10",
"10",
"10",
"01",
"01",
"01",
"10",
"10",
"10",
"00",
"10",
"00",
"01",
"00",
"10",
"11",
"01",
"11",
"01",
"00",
"00",
"00",
"00",
"10",
"11",
"10",
"11",
"10",
"01",
"00",
"00",
"11",
"01",
"10",
"01",
"10",
"00",
"10",
"00",
"01",
"00",
"11",
"10",
"10",
"00",
"10",
"01",
"01",
"11",
"10",
"00",
"10",
"11",
"01",
"01",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"00",
"10",
"11",
"11",
"01",
"11",
"10",
"11",
"11",
"10",
"00",
"00",
"10",
"00",
"11",
"00",
"10",
"00",
"11",
"01",
"10",
"01",
"10",
"11",
"10",
"10",
"00",
"01",
"00",
"11",
"01",
"10",
"01",
"01",
"00",
"10",
"10",
"11",
"10",
"00",
"10",
"11",
"00",
"01",
"01",
"00",
"10",
"11",
"11",
"00",
"11",
"01",
"00",
"11",
"00",
"01",
"11",
"10",
"00",
"11",
"11",
"00",
"00",
"00",
"10",
"10",
"00",
"10",
"00",
"10",
"00",
"00",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"11",
"00",
"11",
"01",
"10",
"00",
"00",
"10",
"10",
"10",
"00",
"01",
"11",
"00",
"00",
"01",
"00",
"10",
"01",
"01",
"00",
"00",
"10",
"11",
"10",
"01",
"11",
"11",
"10",
"01",
"10",
"01",
"00",
"00",
"11",
"11",
"11",
"10",
"11",
"10",
"11",
"10",
"00",
"01",
"01",
"01",
"10",
"01",
"00",
"00",
"11",
"00",
"10",
"01",
"00",
"11",
"00",
"11",
"10",
"10",
"11",
"11",
"10",
"11",
"11",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"01",
"11",
"00",
"00",
"10",
"10",
"10",
"01",
"10",
"01",
"01",
"10",
"10",
"11",
"00",
"01",
"01",
"11",
"11",
"11",
"01",
"01",
"00",
"11",
"00",
"00",
"11",
"01",
"10",
"00",
"00",
"10",
"01",
"11",
"01",
"11",
"11",
"10",
"01",
"11",
"00",
"10",
"11",
"00",
"11",
"01",
"00",
"01",
"00",
"00",
"10",
"11",
"00",
"11",
"11",
"01",
"10",
"01",
"00",
"00",
"10",
"01",
"11",
"11",
"10",
"10",
"10",
"10",
"01",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"01",
"00",
"01",
"10",
"11",
"01",
"01",
"00",
"01",
"10",
"01",
"01",
"10",
"11",
"01",
"10",
"10",
"00",
"10",
"00",
"00",
"00",
"00",
"11",
"10",
"01",
"11",
"00",
"00",
"10",
"01",
"10",
"00",
"11",
"11",
"10",
"10",
"00",
"10",
"01",
"11",
"01",
"10",
"10",
"11",
"00",
"11",
"00",
"00",
"11",
"11",
"00",
"01",
"01",
"01",
"00",
"11",
"10",
"11",
"10",
"11",
"00",
"01",
"11",
"11",
"01",
"00",
"00",
"01",
"01",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"00",
"10",
"11",
"10",
"00",
"01",
"11",
"01",
"00",
"10",
"10",
"01",
"11",
"11",
"00",
"00",
"10",
"11",
"11",
"00",
"11",
"00",
"11",
"00",
"00",
"11",
"11",
"01",
"00",
"10",
"10",
"00",
"11",
"00",
"11",
"00",
"01",
"11",
"01",
"10",
"11",
"10",
"00",
"01",
"11",
"00",
"01",
"01",
"10",
"01",
"00",
"00",
"10",
"00",
"01",
"01",
"00",
"01",
"00",
"11",
"11",
"11",
"00",
"11",
"00",
"10",
"10",
"10",
"11",
"00",
"10",
"01",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"10",
"11",
"00",
"11",
"10",
"01",
"10",
"10",
"00",
"01",
"00",
"01",
"01",
"11",
"01",
"11",
"00",
"11",
"10",
"01",
"11",
"00",
"10",
"01",
"00",
"11",
"10",
"01",
"10",
"11",
"10",
"01",
"00",
"10",
"10",
"11",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"10",
"11",
"10",
"11",
"01",
"00",
"10",
"01",
"11",
"10",
"11",
"10",
"11",
"11",
"11",
"00",
"11",
"00",
"01",
"01",
"10",
"01",
"00",
"11",
"00",
"10",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"00",
"00",
"10",
"10",
"00",
"11",
"00",
"10",
"00",
"01",
"11",
"00",
"00",
"11",
"10",
"00",
"00",
"01",
"10",
"00",
"01",
"11",
"11",
"11",
"00",
"00",
"11",
"01",
"00",
"01",
"00",
"10",
"10",
"10",
"00",
"01",
"11",
"11",
"01",
"10",
"00",
"01",
"00",
"11",
"01",
"10",
"11",
"11",
"00",
"11",
"01",
"11",
"10",
"11",
"10",
"00",
"11",
"10",
"11",
"00",
"00",
"00",
"00",
"11",
"11",
"00",
"11",
"00",
"10",
"11",
"00",
"01",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"10",
"11",
"00",
"00",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"01",
"11",
"00",
"00",
"00",
"11",
"11",
"10",
"00",
"00",
"11",
"10",
"11",
"11",
"00",
"10",
"00",
"01",
"00",
"01",
"00",
"00",
"00",
"11",
"10",
"01",
"11",
"01",
"00",
"10",
"01",
"11",
"00",
"10",
"01",
"10",
"11",
"10",
"10",
"10",
"00",
"11",
"01",
"11",
"00",
"01",
"10",
"10",
"01",
"11",
"11",
"00",
"11",
"11",
"00",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"10",
"00",
"00",
"10",
"00",
"00",
"11",
"01",
"10",
"00",
"00",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"11",
"11",
"01",
"10",
"11",
"00",
"01",
"00",
"11",
"01",
"01",
"10",
"00",
"00",
"01",
"00",
"01",
"00",
"11",
"11",
"10",
"00",
"11",
"11",
"00",
"00",
"11",
"11",
"00",
"10",
"00",
"01",
"00",
"01",
"00",
"11",
"01",
"10",
"00",
"10",
"10",
"11",
"10",
"00",
"01",
"11",
"10",
"01",
"10",
"01",
"10",
"10",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"10",
"01",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"01",
"10",
"01",
"00",
"11",
"00",
"01",
"00",
"10",
"01",
"11",
"10",
"10",
"11",
"11",
"01",
"00",
"11",
"11",
"01",
"10",
"11",
"00",
"10",
"00",
"11",
"00",
"10",
"10",
"10",
"00",
"11",
"11",
"10",
"00",
"11",
"00",
"10",
"11",
"01",
"01",
"00",
"00",
"11",
"10",
"01",
"10",
"00",
"00",
"01",
"11",
"01",
"10",
"00",
"01",
"10",
"11",
"10",
"10",
"11",
"01",
"00",
"00",
"00",
"10",
"10",
"10",
"01",
"11",
"00",
"01",
"01",
"01",
"00",
"00",
"00",
"11",
"00",
"11",
"00",
"11",
"10",
"11",
"00",
"11",
"01",
"01",
"10",
"00",
"11",
"01",
"10",
"01",
"00",
"10",
"11",
"11",
"01",
"00",
"11",
"10",
"10",
"10",
"10",
"10",
"01",
"00",
"01",
"10",
"11",
"01",
"00",
"01",
"00",
"10",
"11",
"01",
"01",
"00",
"10",
"01",
"01",
"00",
"00",
"10",
"10",
"01",
"10",
"10",
"10",
"11",
"11",
"10",
"00",
"00",
"11",
"01",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"00",
"11",
"00",
"00",
"11",
"10",
"01",
"01",
"01",
"00",
"00",
"01",
"11",
"10",
"10",
"01",
"00",
"10",
"00",
"01",
"11",
"11",
"01",
"10",
"00",
"11",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"10",
"10",
"01",
"10",
"00",
"00",
"01",
"10",
"10",
"10",
"00",
"01",
"11",
"01",
"01",
"00",
"11",
"00",
"11",
"00",
"11",
"11",
"11",
"00",
"00",
"00",
"11",
"00",
"10",
"10",
"11",
"01",
"01",
"10",
"01",
"11",
"00",
"00",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"11",
"10",
"10",
"10",
"00",
"11",
"01",
"10",
"00",
"11",
"01",
"00",
"10",
"11",
"01",
"01",
"10",
"11",
"01",
"00",
"11",
"10",
"10",
"00",
"11",
"00",
"11",
"11",
"11",
"10",
"00",
"01",
"01",
"00",
"00",
"11",
"11",
"11",
"11",
"01",
"11",
"10",
"11",
"00",
"10",
"01",
"01",
"11",
"00",
"10",
"00",
"00",
"10",
"00",
"00",
"01",
"10",
"10",
"01",
"11",
"11",
"11",
"10",
"01",
"00",
"10",
"10",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"11",
"01",
"00",
"11",
"01",
"01",
"00",
"00",
"00",
"11",
"00",
"10",
"00",
"11",
"00",
"00",
"10",
"11",
"11",
"10",
"01",
"10",
"01",
"00",
"00",
"10",
"00",
"11",
"01",
"00",
"10",
"00",
"11",
"01",
"01",
"11",
"01",
"01",
"10",
"10",
"00",
"11",
"10",
"01",
"00",
"10",
"01",
"10",
"01",
"10",
"00",
"00",
"10",
"11",
"01",
"10",
"01",
"10",
"10",
"01",
"11",
"01",
"10",
"10",
"00",
"10",
"01",
"01",
"00",
"11",
"11",
"00",
"11",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"01",
"10",
"11",
"10",
"11",
"00",
"11",
"11",
"11",
"00",
"10",
"11",
"10",
"10",
"11",
"01",
"00",
"11",
"10",
"10",
"10",
"10",
"10",
"11",
"01",
"01",
"01",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"10",
"01",
"00",
"11",
"11",
"10",
"01",
"00",
"10",
"01",
"01",
"11",
"11",
"00",
"11",
"01",
"00",
"01",
"11",
"01",
"10",
"01",
"01",
"11",
"00",
"01",
"01",
"10",
"11",
"00",
"00",
"11",
"11",
"00",
"11",
"01",
"00",
"00",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"00",
"00",
"11",
"00",
"01",
"00",
"10",
"00",
"10",
"00",
"11",
"10",
"10",
"11",
"10",
"00",
"11",
"00",
"10",
"00",
"00",
"11",
"01",
"10",
"00",
"00",
"10",
"10",
"10",
"01",
"11",
"11",
"01",
"01",
"10",
"10",
"10",
"11",
"10",
"01",
"11",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"01",
"00",
"11",
"00",
"10",
"01",
"11",
"11",
"00",
"10",
"00",
"00",
"11",
"01",
"00",
"01",
"01",
"01",
"10",
"11",
"11",
"01",
"01",
"01",
"00",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"10",
"01",
"00",
"10",
"11",
"10",
"10",
"00",
"11",
"11",
"01",
"11",
"11",
"01",
"11",
"00",
"10",
"11",
"10",
"10",
"00",
"11",
"10",
"11",
"11",
"01",
"10",
"10",
"10",
"11",
"00",
"00",
"10",
"10",
"10",
"11",
"01",
"01",
"10",
"10",
"00",
"01",
"01",
"00",
"00",
"10",
"01",
"11",
"10",
"10",
"01",
"00",
"00",
"10",
"10",
"10",
"00",
"11",
"01",
"01",
"00",
"01",
"11",
"10",
"10",
"11",
"10",
"10",
"11",
"11",
"01",
"01",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"00",
"10",
"11",
"00",
"10",
"10",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"10",
"10",
"11",
"10",
"01",
"11",
"11",
"11",
"10",
"11",
"11",
"10",
"11",
"11",
"01",
"10",
"11",
"10",
"01",
"01",
"10",
"00",
"00",
"00",
"01",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"01",
"10",
"01",
"00",
"11",
"10",
"10",
"00",
"10",
"11",
"10",
"01",
"11",
"11",
"01",
"10",
"11",
"10",
"10",
"10",
"11",
"10",
"01",
"10",
"00",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"11",
"11",
"10",
"01",
"00",
"01",
"00",
"01",
"01",
"11",
"11",
"10",
"01",
"00",
"11",
"10",
"01",
"01",
"00",
"11",
"11",
"11",
"11",
"01",
"11",
"00",
"01",
"10",
"00",
"00",
"10",
"01",
"10",
"11",
"01",
"01",
"00",
"10",
"10",
"11",
"01",
"01",
"10",
"01",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"10",
"10",
"10",
"00",
"11",
"00",
"00",
"10",
"11",
"00",
"00",
"01",
"10",
"11",
"11",
"11",
"00",
"00",
"10",
"11",
"10",
"11",
"00",
"11",
"00",
"00",
"01",
"01",
"01",
"10",
"10",
"00",
"00",
"10",
"01",
"10",
"10",
"01",
"11",
"10",
"00",
"01",
"10",
"11",
"01",
"10",
"11",
"10",
"00",
"11",
"11",
"10",
"11",
"11",
"00",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"00",
"11",
"11",
"00",
"00",
"11",
"11",
"10",
"11",
"10",
"11",
"01",
"10",
"11",
"10",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"00",
"10",
"11",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"01",
"11",
"11",
"00",
"01",
"01",
"10",
"01",
"10",
"10",
"01",
"00",
"00",
"00",
"01",
"00",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"01",
"01",
"01",
"01",
"10",
"10",
"01",
"11",
"00",
"01",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"11",
"01",
"00",
"01",
"10",
"11",
"10",
"10",
"01",
"01",
"00",
"01",
"10",
"00",
"10",
"01",
"10",
"11",
"00",
"11",
"01",
"00",
"10",
"11",
"11",
"11",
"11",
"10",
"01",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"01",
"00",
"00",
"10",
"01",
"01",
"11",
"11",
"11",
"00",
"00",
"00",
"00",
"01",
"00",
"00",
"01",
"10",
"10",
"10",
"10",
"00",
"10",
"01",
"00",
"11",
"01",
"00",
"00",
"10",
"01",
"01",
"10",
"10",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"01",
"10",
"11",
"11",
"10",
"00",
"11",
"10",
"00",
"01",
"10",
"01",
"10",
"10",
"00",
"01",
"10",
"00",
"10",
"00",
"00",
"10",
"11",
"10",
"01",
"00",
"10",
"00",
"01",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"11",
"00",
"01",
"00",
"00",
"00",
"00",
"11",
"00",
"01",
"01",
"00",
"00",
"01",
"10",
"00",
"11",
"10",
"01",
"11",
"11",
"11",
"10",
"10",
"11",
"11",
"01",
"00",
"01",
"00",
"00",
"01",
"00",
"00",
"00",
"10",
"11",
"10",
"01",
"00",
"00",
"01",
"10",
"00",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"00",
"11",
"00",
"01",
"11",
"00",
"11",
"01",
"10",
"01",
"01",
"11",
"11",
"11",
"11",
"11",
"10",
"00",
"11",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"10",
"00",
"11",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"01",
"01",
"10",
"11",
"00",
"11",
"00",
"10",
"11",
"11",
"10",
"00",
"11",
"10",
"10",
"11",
"00",
"00",
"10",
"01",
"00",
"10",
"00",
"01",
"11",
"11",
"10",
"01",
"00",
"10",
"10",
"11",
"00",
"11",
"10",
"01",
"01",
"11",
"00",
"11",
"00",
"01",
"11",
"11",
"01",
"00",
"11",
"00",
"00",
"01",
"11",
"10",
"00",
"00",
"01",
"11",
"11",
"11",
"11",
"11",
"01",
"01",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"10",
"01",
"00",
"11",
"11",
"00",
"00",
"01",
"01",
"10",
"01",
"10",
"01",
"11",
"00",
"10",
"00",
"01",
"11",
"00",
"10",
"01",
"10",
"00",
"01",
"10",
"10",
"00",
"10",
"10",
"00",
"11",
"00",
"10",
"01",
"11",
"11",
"01",
"01",
"10",
"11",
"11",
"00",
"00",
"00",
"10",
"01",
"00",
"01",
"10",
"11",
"11",
"01",
"11",
"11",
"00",
"00",
"10",
"11",
"01",
"11",
"10",
"01",
"11",
"11",
"10",
"10",
"11",
"10",
"10",
"10",
"00",
"01",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"00",
"10",
"00",
"11",
"11",
"01",
"00",
"10",
"01",
"01",
"01",
"10",
"10",
"01",
"10",
"10",
"10",
"11",
"10",
"00",
"11",
"10",
"11",
"10",
"11",
"00",
"11",
"00",
"11",
"10",
"00",
"01",
"00",
"01",
"01",
"11",
"10",
"01",
"00",
"10",
"10",
"00",
"10",
"00",
"00",
"11",
"11",
"00",
"11",
"11",
"00",
"11",
"11",
"11",
"11",
"00",
"11",
"00",
"11",
"00",
"00",
"11",
"01",
"00",
"10",
"01",
"10",
"10",
"11",
"10",
"01",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"10",
"10",
"00",
"00",
"10",
"10",
"01",
"00",
"10",
"00",
"01",
"00",
"11",
"10",
"10",
"00",
"01",
"11",
"11",
"11",
"00",
"10",
"00",
"11",
"00",
"01",
"01",
"10",
"01",
"10",
"00",
"11",
"10",
"01",
"01",
"00",
"10",
"10",
"10",
"01",
"00",
"11",
"00",
"10",
"00",
"00",
"01",
"00",
"00",
"10",
"10",
"10",
"00",
"01",
"01",
"01",
"00",
"01",
"11",
"01",
"01",
"10",
"11",
"00",
"11",
"11",
"11",
"10",
"10",
"01",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"10",
"01",
"00",
"00",
"01",
"10",
"00",
"00",
"11",
"10",
"10",
"11",
"00",
"11",
"00",
"00",
"00",
"10",
"11",
"00",
"10",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"00",
"11",
"00",
"00",
"10",
"01",
"00",
"00",
"11",
"01",
"01",
"01",
"00",
"11",
"00",
"11",
"10",
"01",
"00",
"11",
"10",
"11",
"00",
"01",
"11",
"01",
"01",
"11",
"01",
"11",
"11",
"01",
"01",
"01",
"00",
"10",
"10",
"11",
"11",
"11",
"00",
"10",
"00",
"11",
"00",
"11",
"11",
"10",
"10",
"10",
"10",
"00",
"01",
"10",
"11",
"00",
"10",
"11",
"00",
"10",
"00",
"10",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"11",
"11",
"11",
"00",
"01",
"01",
"10",
"11",
"00",
"00",
"11",
"00",
"11",
"10",
"11",
"11",
"11",
"10",
"01",
"10",
"00",
"10",
"11",
"10",
"00",
"00",
"01",
"10",
"00",
"11",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"00",
"00",
"11",
"00",
"10",
"11",
"00",
"10",
"11",
"11",
"01",
"10",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"10",
"00",
"01",
"01",
"00",
"00",
"10",
"00",
"11",
"10",
"11",
"01",
"01",
"11",
"10",
"11",
"01",
"00",
"01",
"01",
"01",
"10",
"11",
"11",
"00",
"01",
"10",
"00",
"11",
"00",
"00",
"11",
"00",
"11",
"01",
"10",
"11",
"00",
"01",
"10",
"11",
"01",
"10",
"11",
"11",
"01",
"11",
"11",
"10",
"10",
"00",
"00",
"01",
"10",
"10",
"01",
"01",
"01",
"00",
"00",
"00",
"01",
"10",
"10",
"10",
"00",
"10",
"01",
"11",
"11",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"00",
"00",
"11",
"01",
"01",
"11",
"00",
"10",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"00",
"11",
"01",
"10",
"01",
"00",
"11",
"00",
"00",
"10",
"00",
"10",
"11",
"10",
"00",
"10",
"01",
"10",
"10",
"00",
"11",
"11",
"10",
"01",
"10",
"11",
"01",
"01",
"10",
"11",
"01",
"01",
"00",
"01",
"10",
"11",
"10",
"01",
"10",
"11",
"01",
"11",
"11",
"01",
"00",
"01",
"10",
"10",
"11",
"10",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"11",
"10",
"01",
"00",
"00",
"10",
"01",
"00",
"11",
"10",
"00",
"10",
"11",
"10",
"00",
"11",
"01",
"11",
"11",
"10",
"01",
"01",
"00",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"01",
"11",
"00",
"00",
"10",
"11",
"00",
"10",
"11",
"11",
"01",
"01",
"01",
"10",
"01",
"11",
"00",
"01",
"11",
"01",
"00",
"00",
"10",
"11",
"11",
"10",
"00",
"10",
"11",
"11",
"00",
"10",
"00",
"11",
"01",
"11",
"11",
"01",
"10",
"00",
"10",
"00",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"10",
"10",
"10",
"10",
"11",
"00",
"10",
"01",
"10",
"01",
"00",
"00",
"10",
"10",
"10",
"00",
"11",
"01",
"10",
"11",
"11",
"11",
"10",
"00",
"00",
"10",
"01",
"00",
"00",
"11",
"10",
"01",
"10",
"10",
"01",
"01",
"01",
"01",
"01",
"10",
"10",
"01",
"00",
"11",
"11",
"01",
"10",
"10",
"11",
"01",
"01",
"00",
"11",
"10",
"11",
"00",
"11",
"11",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"01",
"10",
"01",
"10",
"10",
"10",
"00",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"10",
"11",
"10",
"01",
"00",
"00",
"00",
"01",
"11",
"11",
"00",
"01",
"01",
"11",
"11",
"00",
"01",
"01",
"01",
"01",
"10",
"01",
"10",
"01",
"10",
"11",
"11",
"00",
"10",
"01",
"10",
"10",
"11",
"11",
"10",
"10",
"01",
"01",
"00",
"01",
"11",
"10",
"00",
"01",
"00",
"01",
"10",
"00",
"01",
"10",
"10",
"10",
"10",
"11",
"10",
"11",
"00",
"10",
"01",
"11",
"10",
"00",
"01",
"01",
"11",
"10",
"11",
"01",
"11",
"11",
"01",
"11",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"10",
"11",
"00",
"10",
"01",
"01",
"11",
"01",
"10",
"00",
"00",
"00",
"10",
"10",
"00",
"10",
"01",
"11",
"00",
"11",
"11",
"11",
"00",
"10",
"10",
"00",
"01",
"11",
"00",
"10",
"00",
"01",
"00",
"11",
"11",
"01",
"00",
"11",
"00",
"00",
"01",
"01",
"00",
"11",
"10",
"00",
"10",
"10",
"00",
"10",
"01",
"11",
"10",
"10",
"00",
"01",
"11",
"11",
"01",
"01",
"01",
"01",
"10",
"00",
"01",
"11",
"10",
"01",
"11",
"10",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"11",
"00",
"11",
"11",
"10",
"10",
"10",
"11",
"01",
"11",
"11",
"01",
"10",
"10",
"01",
"01",
"00",
"00",
"01",
"10",
"00",
"01",
"00",
"11",
"10",
"01",
"11",
"10",
"11",
"01",
"00",
"00",
"01",
"11",
"01",
"00",
"11",
"01",
"01",
"00",
"01",
"00",
"11",
"01",
"10",
"11",
"00",
"11",
"01",
"01",
"01",
"11",
"11",
"01",
"11",
"01",
"11",
"10",
"10",
"11",
"10",
"11",
"00",
"00",
"10",
"11",
"00",
"11",
"10",
"10",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"01",
"10",
"01",
"11",
"01",
"10",
"11",
"11",
"01",
"01",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"10",
"01",
"00",
"00",
"00",
"00",
"11",
"00",
"11",
"11",
"11",
"11",
"00",
"00",
"00",
"11",
"10",
"11",
"00",
"10",
"01",
"01",
"00",
"11",
"00",
"00",
"11",
"01",
"10",
"00",
"01",
"00",
"11",
"00",
"00",
"01",
"01",
"11",
"00",
"11",
"00",
"10",
"11",
"01",
"10",
"01",
"10",
"11",
"10",
"01",
"11",
"10",
"11",
"00",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"10",
"11",
"11",
"01",
"00",
"01",
"01",
"11",
"00",
"01",
"00",
"00",
"01",
"11",
"11",
"10",
"10",
"01",
"10",
"10",
"01",
"10",
"11",
"01",
"01",
"01",
"00",
"11",
"10",
"10",
"11",
"11",
"10",
"10",
"11",
"00",
"00",
"11",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"11",
"10",
"10",
"10",
"01",
"00",
"01",
"01",
"00",
"11",
"00",
"01",
"11",
"00",
"01",
"10",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"10",
"10",
"10",
"00",
"00",
"10",
"11",
"01",
"01",
"01",
"11",
"01",
"11",
"01",
"11",
"01",
"10",
"01",
"01",
"00",
"01",
"10",
"01",
"00",
"01",
"01",
"11",
"01",
"11",
"10",
"10",
"00",
"00",
"10",
"01",
"01",
"10",
"01",
"00",
"00",
"01",
"00",
"01",
"00",
"00",
"00",
"11",
"10",
"01",
"10",
"11",
"11",
"10",
"10",
"00",
"01",
"00",
"00",
"11",
"00",
"00",
"00",
"10",
"11",
"01",
"10",
"10",
"10",
"10",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"01",
"00",
"00",
"01",
"00",
"11",
"01",
"01",
"11",
"00",
"00",
"00",
"11",
"11",
"11",
"01",
"11",
"00",
"11",
"01",
"11",
"01",
"11",
"10",
"11",
"10",
"10",
"11",
"11",
"10",
"11",
"10",
"00",
"01",
"00",
"11",
"10",
"00",
"01",
"01",
"01",
"10",
"11",
"10",
"11",
"10",
"11",
"00",
"10",
"10",
"11",
"00",
"10",
"11",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"00",
"11",
"01",
"11",
"10",
"01",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"01",
"10",
"11",
"11",
"01",
"01",
"11",
"11",
"00",
"01",
"01",
"00",
"01",
"01",
"11",
"00",
"11",
"01",
"00",
"11",
"01",
"11",
"01",
"11",
"10",
"00",
"01",
"11",
"01",
"10",
"10",
"01",
"11",
"01",
"00",
"00",
"01",
"11",
"00",
"10",
"00",
"01",
"01",
"00",
"11",
"11",
"01",
"00",
"00",
"11",
"01",
"10",
"11",
"11",
"00",
"11",
"01",
"00",
"01",
"01",
"10",
"10",
"11",
"10",
"10",
"00",
"01",
"01",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"10",
"00",
"00",
"11",
"01",
"11",
"11",
"00",
"11",
"00",
"10",
"01",
"11",
"00",
"00",
"01",
"11",
"01",
"01",
"10",
"01",
"01",
"10",
"10",
"10",
"01",
"10",
"00",
"11",
"00",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"11",
"10",
"00",
"10",
"01",
"01",
"10",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"10",
"00",
"10",
"11",
"11",
"00",
"11",
"10",
"01",
"10",
"00",
"00",
"11",
"10",
"01",
"11",
"01",
"00",
"10",
"10",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"01",
"11",
"00",
"01",
"01",
"11",
"00",
"10",
"01",
"11",
"00",
"11",
"00",
"01",
"01",
"00",
"10",
"11",
"10",
"11",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"01",
"11",
"11",
"11",
"00",
"00",
"01",
"00",
"11",
"10",
"10",
"11",
"01",
"00",
"10",
"10",
"11",
"00",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"11",
"10",
"11",
"10",
"10",
"01",
"01",
"10",
"10",
"00",
"10",
"11",
"10",
"11",
"01",
"10",
"01",
"10",
"01",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"00",
"00",
"10",
"00",
"01",
"11",
"00",
"10",
"11",
"11",
"10",
"11",
"01",
"00",
"00",
"01",
"11",
"10",
"00",
"00",
"11",
"10",
"01",
"11",
"00",
"00",
"01",
"11",
"10",
"11",
"10",
"10",
"01",
"11",
"01",
"01",
"11",
"11",
"00",
"00",
"10",
"11",
"11",
"10",
"01",
"10",
"11",
"10",
"10",
"11",
"10",
"01",
"10",
"00",
"10",
"00",
"00",
"00",
"11",
"11",
"11",
"11",
"00",
"01",
"11",
"00",
"01",
"00",
"10",
"01",
"01",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"01",
"01",
"01",
"10",
"01",
"11",
"11",
"10",
"00",
"01",
"01",
"00",
"11",
"10",
"11",
"10",
"00",
"01",
"00",
"01",
"10",
"00",
"11",
"01",
"01",
"00",
"11",
"11",
"10",
"11",
"01",
"00",
"01",
"11",
"11",
"00",
"00",
"01",
"01",
"01",
"11",
"00",
"00",
"11",
"01",
"10",
"10",
"10",
"00",
"01",
"01",
"11",
"10",
"01",
"10",
"01",
"01",
"00",
"10",
"00",
"11",
"10",
"00",
"10",
"10",
"01",
"01",
"00",
"01",
"00",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"10",
"00",
"01",
"00",
"10",
"00",
"10",
"00",
"10",
"11",
"11",
"01",
"00",
"00",
"10",
"10",
"11",
"10",
"00",
"00",
"10",
"01",
"11",
"11",
"01",
"11",
"00",
"00",
"11",
"01",
"11",
"01",
"00",
"00",
"10",
"10",
"00",
"00",
"10",
"10",
"00",
"00",
"00",
"00",
"10",
"00",
"01",
"10",
"00",
"00",
"11",
"00",
"00",
"11",
"11",
"00",
"10",
"11",
"01",
"01",
"01",
"01",
"11",
"00",
"11",
"10",
"10",
"10",
"11",
"01",
"00",
"00",
"01",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"10",
"11",
"11",
"00",
"00",
"10",
"00",
"00",
"01",
"01",
"00",
"10",
"01",
"11",
"00",
"11",
"01",
"00",
"01",
"00",
"00",
"01",
"10",
"01",
"00",
"01",
"01",
"10",
"11",
"10",
"00",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"00",
"00",
"11",
"10",
"11",
"00",
"01",
"00",
"10",
"00",
"11",
"10",
"10",
"11",
"00",
"00",
"11",
"10",
"11",
"00",
"11",
"10",
"00",
"00",
"10",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"10",
"00",
"00",
"10",
"00",
"01",
"11",
"10",
"01",
"11",
"10",
"01",
"10",
"01",
"10",
"01",
"00",
"01",
"11",
"10",
"11",
"01",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"00",
"10",
"11",
"00",
"00",
"10",
"00",
"10",
"10",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"10",
"10",
"01",
"00",
"11",
"11",
"01",
"01",
"00",
"11",
"11",
"10",
"00",
"10",
"00",
"10",
"10",
"00",
"10",
"01",
"11",
"00",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"01",
"00",
"00",
"00",
"01",
"11",
"10",
"00",
"00",
"00",
"11",
"11",
"11",
"01",
"10",
"10",
"11",
"10",
"00",
"11",
"00",
"10",
"11",
"01",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"10",
"10",
"00",
"11",
"11",
"00",
"10",
"00",
"01",
"00",
"01",
"01",
"10",
"10",
"11",
"01",
"10",
"00",
"00",
"11",
"10",
"11",
"10",
"11",
"10",
"10",
"10",
"10",
"00",
"00",
"11",
"10",
"10",
"11",
"11",
"11",
"10",
"11",
"01",
"10",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"01",
"00",
"11",
"01",
"10",
"10",
"00",
"10",
"01",
"10",
"01",
"10",
"11",
"10",
"00",
"10",
"10",
"11",
"10",
"11",
"01",
"00",
"10",
"10",
"10",
"00",
"10",
"00",
"10",
"11",
"00",
"10",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"10",
"11",
"00",
"01",
"00",
"11",
"10",
"00",
"10",
"10",
"00",
"11",
"10",
"00",
"00",
"01",
"00",
"10",
"01",
"10",
"11",
"00",
"00",
"01",
"10",
"10",
"11",
"01",
"11",
"10",
"00",
"10",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"11",
"01",
"00",
"00",
"01",
"11",
"00",
"11",
"00",
"10",
"01",
"01",
"10",
"10",
"00",
"10",
"01",
"11",
"00",
"01",
"11",
"11",
"00",
"10",
"11",
"10",
"10",
"01",
"00",
"10",
"10",
"00",
"00",
"01",
"10",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"10",
"01",
"01",
"10",
"01",
"10",
"10",
"00",
"10",
"00",
"11",
"00",
"10",
"11",
"00",
"10",
"01",
"10",
"01",
"10",
"00",
"11",
"00",
"01",
"10",
"00",
"10",
"01",
"10",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"10",
"11",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"11",
"01",
"00",
"10",
"10",
"01",
"11",
"10",
"00",
"01",
"01",
"00",
"00",
"11",
"11",
"00",
"10",
"01",
"00",
"10",
"01",
"01",
"10",
"11",
"00",
"11",
"11",
"01",
"00",
"11",
"10",
"00",
"11",
"10",
"10",
"10",
"00",
"10",
"10",
"01",
"10",
"10",
"10",
"01",
"00",
"00",
"10",
"01",
"11",
"11",
"00",
"01",
"10",
"00",
"11",
"11",
"11",
"01",
"10",
"01",
"00",
"11",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"00",
"01",
"01",
"00",
"00",
"01",
"00",
"11",
"10",
"10",
"10",
"01",
"00",
"10",
"10",
"10",
"01",
"01",
"11",
"00",
"10",
"11",
"11",
"01",
"11",
"00",
"10",
"10",
"10",
"10",
"11",
"00",
"00",
"11",
"11",
"01",
"00",
"11",
"10",
"11",
"10",
"11",
"01",
"01",
"00",
"01",
"00",
"11",
"00",
"00",
"00",
"00",
"01",
"10",
"11",
"00",
"00",
"00",
"01",
"11",
"11",
"11",
"11",
"10",
"10",
"11",
"11",
"10",
"11",
"11",
"00",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"11",
"11",
"00",
"00",
"11",
"01",
"00",
"10",
"11",
"01",
"00",
"11",
"10",
"10",
"00",
"00",
"10",
"10",
"10",
"01",
"01",
"10",
"01",
"11",
"11",
"00",
"11",
"11",
"10",
"01",
"11",
"01",
"01",
"11",
"01",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"01",
"01",
"01",
"00",
"11",
"01",
"01",
"00",
"11",
"11",
"10",
"01",
"10",
"11",
"01",
"11",
"10",
"11",
"10",
"00",
"10",
"00",
"01",
"01",
"01",
"10",
"10",
"00",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"10",
"11",
"01",
"10",
"11",
"11",
"10",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"10",
"00",
"01",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"11",
"01",
"11",
"11",
"10",
"01",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"11",
"00",
"01",
"01",
"00",
"00",
"00",
"11",
"01",
"00",
"10",
"00",
"01",
"01",
"01",
"00",
"11",
"10",
"11",
"00",
"11",
"10",
"10",
"10",
"01",
"10",
"01",
"01",
"01",
"11",
"01",
"11",
"10",
"11",
"01",
"10",
"01",
"11",
"11",
"11",
"11",
"00",
"01",
"01",
"10",
"10",
"00",
"11",
"11",
"11",
"00",
"11",
"11",
"01",
"10",
"11",
"01",
"10",
"10",
"01",
"10",
"00",
"11",
"10",
"00",
"01",
"01",
"11",
"00",
"01",
"10",
"00",
"00",
"01",
"10",
"11",
"00",
"00",
"10",
"10",
"10",
"00",
"01",
"10",
"10",
"11",
"00",
"11",
"01",
"11",
"00",
"10",
"11",
"10",
"10",
"00",
"01",
"11",
"10",
"00",
"10",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"11",
"00",
"10",
"11",
"00",
"01",
"11",
"11",
"11",
"00",
"10",
"00",
"10",
"00",
"11",
"00",
"11",
"00",
"10",
"00",
"00",
"10",
"01",
"00",
"11",
"01",
"11",
"00",
"00",
"11",
"01",
"01",
"01",
"00",
"00",
"01",
"11",
"00",
"11",
"11",
"11",
"01",
"00",
"00",
"01",
"11",
"01",
"11",
"00",
"01",
"00",
"11",
"10",
"00",
"00",
"01",
"11",
"01",
"01",
"00",
"01",
"00",
"00",
"11",
"01",
"10",
"01",
"10",
"01",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"11",
"00",
"10",
"11",
"01",
"01",
"01",
"11",
"00",
"10",
"10",
"01",
"00",
"01",
"11",
"10",
"01",
"00",
"00",
"11",
"01",
"11",
"10",
"10",
"01",
"11",
"01",
"01",
"10",
"00",
"00",
"10",
"01",
"00",
"00",
"10",
"01",
"00",
"00",
"01",
"10",
"11",
"01",
"01",
"11",
"01",
"01",
"01",
"00",
"01",
"10",
"10",
"10",
"00",
"11",
"01",
"00",
"01",
"10",
"10",
"01",
"10",
"10",
"00",
"00",
"10",
"00",
"10",
"00",
"00",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"01",
"11",
"01",
"10",
"11",
"11",
"01",
"10",
"01",
"01",
"10",
"00",
"11",
"11",
"00",
"10",
"00",
"11",
"01",
"10",
"10",
"10",
"10",
"11",
"00",
"01",
"01",
"10",
"00",
"00",
"11",
"10",
"11",
"10",
"01",
"00",
"00",
"10",
"10",
"10",
"11",
"10",
"10",
"01",
"00",
"00",
"10",
"01",
"11",
"00",
"00",
"10",
"10",
"00",
"01",
"11",
"10",
"11",
"10",
"11",
"01",
"00",
"10",
"10",
"10",
"10",
"11",
"10",
"11",
"00",
"00",
"10",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"00",
"01",
"01",
"01",
"00",
"00",
"11",
"11",
"01",
"00",
"10",
"11",
"11",
"11",
"10",
"11",
"00",
"10",
"01",
"00",
"10",
"01",
"10",
"01",
"10",
"00",
"00",
"11",
"01",
"01",
"00",
"01",
"01",
"10",
"10",
"00",
"10",
"00",
"11",
"10",
"11",
"01",
"11",
"01",
"01",
"01",
"01",
"01",
"01",
"00",
"11",
"10",
"00",
"00",
"10",
"01",
"01",
"11",
"10",
"11",
"01",
"10",
"00",
"01",
"11",
"01",
"00",
"01",
"10",
"00",
"01",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"10",
"01",
"00",
"11",
"01",
"00",
"00",
"01",
"01",
"01",
"11",
"11",
"00",
"00",
"01",
"11",
"00",
"01",
"01",
"11",
"10",
"00",
"10",
"00",
"01",
"10",
"11",
"11",
"11",
"11",
"01",
"10",
"01",
"00",
"01",
"11",
"11",
"10",
"10",
"11",
"10",
"10",
"00",
"01",
"10",
"00",
"00",
"11",
"01",
"10",
"00",
"10",
"01",
"10",
"10",
"00",
"01",
"10",
"00",
"10",
"01",
"11",
"01",
"10",
"01",
"10",
"00",
"11",
"00",
"11",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"00",
"01",
"00",
"00",
"11",
"10",
"01",
"10",
"10",
"10",
"00",
"00",
"10",
"11",
"10",
"10",
"10",
"01",
"11",
"00",
"00",
"01",
"01",
"01",
"11",
"11",
"01",
"11",
"01",
"11",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"00",
"11",
"01",
"01",
"01",
"10",
"00",
"11",
"00",
"01",
"11",
"00",
"01",
"10",
"10",
"00",
"10",
"01",
"00",
"00",
"01",
"11",
"00",
"10",
"00",
"00",
"00",
"01",
"00",
"10",
"00",
"10",
"10",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"01",
"00",
"11",
"01",
"00",
"01",
"10",
"11",
"10",
"10",
"01",
"10",
"01",
"10",
"11",
"00",
"00",
"01",
"10",
"11",
"11",
"00",
"00",
"10",
"10",
"00",
"11",
"01",
"11",
"11",
"01",
"00",
"10",
"11",
"01",
"00",
"00",
"10",
"10",
"10",
"10",
"01",
"00",
"10",
"01",
"10",
"11",
"11",
"10",
"11",
"00",
"10",
"10",
"01",
"00",
"01",
"11",
"11",
"01",
"11",
"11",
"01",
"00",
"10",
"11",
"00",
"10",
"10",
"11",
"00",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"11",
"10",
"00",
"00",
"01",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"10",
"11",
"01",
"11",
"01",
"10",
"10",
"10",
"11",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"11",
"00",
"01",
"11",
"01",
"01",
"11",
"01",
"01",
"10",
"10",
"11",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"10",
"00",
"01",
"01",
"01",
"01",
"00",
"00",
"01",
"00",
"10",
"01",
"00",
"01",
"10",
"00",
"11",
"00",
"11",
"00",
"10",
"10",
"11",
"10",
"00",
"01",
"00",
"00",
"01",
"00",
"00",
"01",
"00",
"00",
"10",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"10",
"00",
"00",
"10",
"10",
"11",
"11",
"10",
"00",
"11",
"01",
"11",
"00",
"10",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"00",
"10",
"11",
"01",
"00",
"11",
"01",
"11",
"11",
"00",
"01",
"10",
"00",
"01",
"00",
"00",
"01",
"10",
"00",
"11",
"01",
"10",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"10",
"10",
"10",
"10",
"01",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"10",
"01",
"10",
"00",
"11",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"00",
"10",
"00",
"01",
"11",
"01",
"01",
"00",
"01",
"10",
"11",
"01",
"00",
"10",
"11",
"10",
"11",
"11",
"01",
"01",
"00",
"01",
"11",
"01",
"10",
"01",
"10",
"11",
"10",
"01",
"00",
"10",
"00",
"01",
"00",
"10",
"11",
"10",
"00",
"01",
"11",
"11",
"11",
"00",
"01",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"00",
"10",
"00",
"00",
"01",
"11",
"10",
"01",
"01",
"11",
"00",
"01",
"11",
"01",
"10",
"00",
"00",
"11",
"01",
"10",
"00",
"10",
"01",
"01",
"01",
"10",
"01",
"11",
"01",
"10",
"11",
"10",
"10",
"00",
"00",
"11",
"00",
"11",
"00",
"10",
"11",
"10",
"11",
"00",
"10",
"10",
"10",
"00",
"00",
"11",
"01",
"01",
"01",
"11",
"11",
"01",
"00",
"00",
"11",
"01",
"01",
"11",
"01",
"00",
"10",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"10",
"01",
"11",
"10",
"01",
"11",
"00",
"11",
"11",
"11",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"11",
"10",
"11",
"00",
"11",
"00",
"01",
"01",
"10",
"01",
"10",
"10",
"01",
"00",
"11",
"00",
"00",
"01",
"10",
"10",
"11",
"00",
"01",
"11",
"10",
"10",
"01",
"10",
"00",
"01",
"01",
"00",
"01",
"01",
"11",
"01",
"11",
"11",
"00",
"01",
"10",
"10",
"00",
"00",
"11",
"10",
"01",
"11",
"01",
"00",
"01",
"10",
"01",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"01",
"00",
"00",
"00",
"01",
"01",
"11",
"01",
"11",
"11",
"11",
"01",
"11",
"00",
"00",
"11",
"00",
"01",
"01",
"01",
"11",
"01",
"11",
"10",
"01",
"11",
"00",
"00",
"00",
"00",
"10",
"00",
"00",
"10",
"01",
"00",
"11",
"11",
"11",
"01",
"01",
"11",
"01",
"00",
"10",
"10",
"00",
"11",
"01",
"01",
"10",
"01",
"10",
"10",
"00",
"10",
"11",
"11",
"00",
"11",
"10",
"11",
"00",
"11",
"00",
"00",
"00",
"11",
"00",
"01",
"01",
"11",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"10",
"11",
"01",
"00",
"01",
"10",
"11",
"00",
"01",
"01",
"00",
"10",
"00",
"00",
"10",
"10",
"11",
"11",
"01",
"01",
"11",
"00",
"11",
"10",
"11",
"10",
"11",
"10",
"10",
"01",
"11",
"01",
"10",
"11",
"11",
"00",
"10",
"11",
"01",
"00",
"00",
"10",
"10",
"00",
"01",
"01",
"11",
"10",
"10",
"00",
"10",
"10",
"00",
"01",
"11",
"11",
"01",
"01",
"00",
"10",
"10",
"01",
"10",
"11",
"00",
"01",
"01",
"01",
"10",
"10",
"00",
"00",
"10",
"01",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"01",
"11",
"10",
"10",
"10",
"11",
"01",
"00",
"00",
"01",
"00",
"00",
"00",
"01",
"11",
"01",
"00",
"00",
"00",
"01",
"01",
"10",
"00",
"11",
"10",
"00",
"10",
"01",
"11",
"01",
"00",
"11",
"10",
"11",
"11",
"01",
"10",
"10",
"11",
"01",
"00",
"11",
"11",
"10",
"10",
"01",
"00",
"01",
"01",
"10",
"10",
"10",
"11",
"01",
"00",
"11",
"00",
"01",
"00",
"10",
"11",
"10",
"00",
"01",
"10",
"01",
"11",
"11",
"01",
"01",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"00",
"10",
"01",
"00",
"00",
"10",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"00",
"10",
"11",
"00",
"01",
"00",
"00",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"01",
"10",
"01",
"11",
"00",
"10",
"01",
"00",
"00",
"11",
"10",
"10",
"01",
"00",
"10",
"00",
"11",
"01",
"10",
"11",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"10",
"10",
"00",
"11",
"10",
"00",
"10",
"10",
"11",
"00",
"00",
"01",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"00",
"01",
"01",
"10",
"11",
"10",
"00",
"10",
"01",
"11",
"10",
"10",
"00",
"00",
"00",
"11",
"01",
"10",
"00",
"11",
"10",
"00",
"01",
"01",
"10",
"01",
"10",
"01",
"10",
"00",
"11",
"00",
"10",
"00",
"01",
"01",
"01",
"10",
"11",
"10",
"11",
"11",
"10",
"00",
"11",
"00",
"10",
"00",
"11",
"00",
"00",
"11",
"10",
"11",
"10",
"10",
"01",
"01",
"11",
"10",
"10",
"10",
"11",
"01",
"01",
"01",
"11",
"10",
"00",
"11",
"01",
"01",
"10",
"10",
"10",
"11",
"00",
"01",
"01",
"11",
"01",
"10",
"11",
"10",
"11",
"00",
"00",
"01",
"00",
"11",
"00",
"10",
"00",
"00",
"11",
"11",
"00",
"01",
"11",
"00",
"10",
"00",
"00",
"01",
"10",
"01",
"11",
"10",
"00",
"00",
"11",
"00",
"01",
"01",
"10",
"11",
"10",
"11",
"00",
"00",
"10",
"00",
"11",
"11",
"10",
"00",
"10",
"11",
"00",
"11",
"10",
"01",
"10",
"00",
"00",
"11",
"11",
"01",
"01",
"00",
"10",
"11",
"01",
"11",
"11",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"10",
"00",
"00",
"00",
"10",
"00",
"10",
"01",
"00",
"01",
"00",
"11",
"11",
"01",
"01",
"11",
"01",
"01",
"10",
"11",
"00",
"10",
"10",
"00",
"10",
"11",
"00",
"01",
"00",
"10",
"01",
"10",
"11",
"10",
"10",
"00",
"00",
"11",
"11",
"01",
"11",
"10",
"01",
"11",
"10",
"11",
"10",
"00",
"10",
"01",
"01",
"10",
"01",
"01",
"00",
"01",
"10",
"00",
"11",
"00",
"00",
"10",
"01",
"11",
"11",
"11",
"01",
"00",
"11",
"10",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"01",
"00",
"11",
"11",
"10",
"11",
"10",
"01",
"11",
"11",
"10",
"01",
"11",
"11",
"01",
"10",
"01",
"01",
"00",
"01",
"11",
"11",
"00",
"11",
"10",
"01",
"10",
"01",
"00",
"01",
"00",
"10",
"00",
"01",
"01",
"00",
"00",
"00",
"01",
"00",
"10",
"01",
"01",
"00",
"01",
"01",
"11",
"01",
"11",
"10",
"01",
"00",
"00",
"11",
"11",
"10",
"00",
"10",
"11",
"10",
"11",
"10",
"11",
"10",
"01",
"10",
"10",
"10",
"11",
"11",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"01",
"00",
"00",
"10",
"11",
"01",
"10",
"11",
"00",
"01",
"00",
"11",
"01",
"01",
"00",
"11",
"00",
"01",
"11",
"00",
"01",
"00",
"01",
"10",
"11",
"11",
"01",
"10",
"11",
"00",
"01",
"01",
"10",
"01",
"01",
"10",
"11",
"10",
"01",
"10",
"11",
"01",
"11",
"11",
"01",
"11",
"11",
"00",
"11",
"10",
"00",
"10",
"11",
"10",
"00",
"00",
"10",
"00",
"10",
"11",
"00",
"10",
"01",
"11",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"11",
"10",
"00",
"00",
"01",
"01",
"01",
"00",
"01",
"10",
"00",
"00",
"01",
"01",
"00",
"00",
"00",
"10",
"10",
"01",
"10",
"11",
"10",
"11",
"11",
"00",
"10",
"00",
"00",
"10",
"10",
"00",
"10",
"11",
"10",
"00",
"11",
"10",
"11",
"01",
"11",
"11",
"10",
"01",
"10",
"11",
"11",
"01",
"10",
"01",
"01",
"00",
"10",
"11",
"00",
"00",
"01",
"00",
"00",
"00",
"10",
"11",
"10",
"00",
"01",
"11",
"10",
"10",
"01",
"00",
"11",
"01",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"00",
"01",
"11",
"10",
"00",
"00",
"00",
"11",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"11",
"01",
"01",
"01",
"11",
"10",
"10",
"00",
"11",
"01",
"11",
"10",
"01",
"01",
"00",
"10",
"01",
"01",
"11",
"00",
"11",
"11",
"10",
"10",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"10",
"10",
"01",
"10",
"11",
"10",
"01",
"01",
"00",
"11",
"00",
"00",
"10",
"00",
"11",
"01",
"11",
"00",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"11",
"10",
"00",
"01",
"10",
"10",
"11",
"11",
"00",
"01",
"11",
"01",
"00",
"10",
"01",
"00",
"11",
"01",
"01",
"00",
"11",
"11",
"10",
"00",
"11",
"00",
"11",
"11",
"00",
"10",
"00",
"11",
"11",
"00",
"01",
"11",
"10",
"01",
"01",
"10",
"10",
"00",
"11",
"11",
"00",
"00",
"01",
"10",
"11",
"10",
"11",
"00",
"00",
"10",
"11",
"00",
"11",
"11",
"11",
"10",
"11",
"01",
"01",
"01",
"00",
"11",
"10",
"11",
"11",
"01",
"10",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"11",
"00",
"00",
"01",
"01",
"10",
"00",
"11",
"00",
"11",
"01",
"00",
"10",
"00",
"01",
"01",
"01",
"01",
"10",
"01",
"10",
"00",
"00",
"01",
"11",
"10",
"00",
"00",
"10",
"10",
"10",
"11",
"01",
"00",
"11",
"00",
"10",
"00",
"10",
"00",
"10",
"00",
"11",
"10",
"01",
"10",
"00",
"00",
"01",
"00",
"11",
"10",
"00",
"10",
"11",
"00",
"01",
"01",
"00",
"01",
"00",
"01",
"00",
"10",
"10",
"11",
"11",
"00",
"11",
"10",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"00",
"00",
"01",
"10",
"01",
"00",
"10",
"00",
"11",
"00",
"11",
"00",
"10",
"00",
"00",
"11",
"10",
"10",
"00",
"10",
"01",
"01",
"10",
"10",
"01",
"00",
"11",
"00",
"10",
"01",
"01",
"11",
"10",
"00",
"01",
"10",
"01",
"11",
"10",
"00",
"10",
"01",
"10",
"01",
"10",
"01",
"10",
"10",
"01",
"00",
"10",
"00",
"00",
"00",
"11",
"01",
"10",
"10",
"10",
"01",
"11",
"01",
"11",
"11",
"01",
"00",
"10",
"00",
"00",
"00",
"10",
"01",
"10",
"11",
"11",
"01",
"10",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"01",
"00",
"00",
"01",
"00",
"01",
"00",
"00",
"01",
"11",
"10",
"11",
"00",
"11",
"01",
"10",
"01",
"00",
"01",
"11",
"10",
"01",
"11",
"01",
"11",
"11",
"01",
"11",
"10",
"10",
"00",
"10",
"11",
"11",
"00",
"11",
"11",
"00",
"00",
"00",
"11",
"10",
"01",
"00",
"10",
"00",
"00",
"00",
"01",
"01",
"00",
"11",
"10",
"01",
"11",
"01",
"01",
"11",
"00",
"11",
"11",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"00",
"00",
"01",
"10",
"01",
"11",
"01",
"11",
"00",
"10",
"01",
"00",
"10",
"11",
"11",
"01",
"00",
"00",
"10",
"10",
"11",
"01",
"01",
"01",
"00",
"10",
"01",
"01",
"00",
"00",
"11",
"11",
"10",
"10",
"10",
"10",
"11",
"11",
"11",
"00",
"10",
"01",
"01",
"10",
"00",
"10",
"11",
"10",
"00",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"11",
"10",
"00",
"01",
"00",
"11",
"10",
"10",
"00",
"00",
"10",
"01",
"01",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"11",
"01",
"00",
"10",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"00",
"01",
"01",
"11",
"01",
"10",
"00",
"01",
"01",
"01",
"11",
"11",
"01",
"00",
"00",
"11",
"00",
"01",
"01",
"11",
"00",
"01",
"01",
"00",
"00",
"01",
"11",
"00",
"10",
"00",
"00",
"10",
"10",
"11",
"00",
"01",
"10",
"01",
"00",
"11",
"01",
"01",
"10",
"11",
"01",
"00",
"10",
"01",
"01",
"00",
"11",
"01",
"11",
"11",
"01",
"11",
"11",
"01",
"11",
"10",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"00",
"11",
"01",
"00",
"10",
"01",
"11",
"00",
"00",
"11",
"10",
"10",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"01",
"01",
"00",
"11",
"00",
"11",
"11",
"01",
"11",
"00",
"10",
"01",
"11",
"10",
"10",
"10",
"01",
"01",
"11",
"11",
"10",
"10",
"10",
"10",
"00",
"00",
"11",
"00",
"00",
"01",
"01",
"10",
"00",
"01",
"00",
"10",
"01",
"01",
"11",
"01",
"10",
"01",
"10",
"11",
"10",
"01",
"01",
"11",
"00",
"00",
"11",
"01",
"10",
"00",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"01",
"10",
"00",
"10",
"00",
"01",
"00",
"00",
"00",
"00",
"11",
"01",
"01",
"11",
"10",
"11",
"11",
"01",
"00",
"11",
"01",
"11",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"10",
"11",
"00",
"10",
"10",
"01",
"00",
"10",
"10",
"10",
"01",
"01",
"10",
"00",
"11",
"00",
"10",
"11",
"11",
"11",
"11",
"01",
"10",
"01",
"00",
"11",
"01",
"10",
"01",
"11",
"11",
"10",
"01",
"01",
"10",
"00",
"01",
"11",
"11",
"10",
"10",
"01",
"10",
"10",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"00",
"10",
"11",
"10",
"10",
"01",
"00",
"10",
"01",
"01",
"01",
"11",
"10",
"10",
"01",
"01",
"10",
"11",
"01",
"01",
"11",
"00",
"00",
"01",
"10",
"00",
"10",
"01",
"01",
"10",
"00",
"10",
"10",
"00",
"11",
"00",
"01",
"01",
"10",
"01",
"00",
"10",
"00",
"00",
"00",
"00",
"10",
"00",
"11",
"10",
"11",
"01",
"11",
"00",
"00",
"10",
"11",
"11",
"10",
"01",
"11",
"11",
"00",
"11",
"10",
"01",
"10",
"00",
"01",
"10",
"11",
"10",
"10",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"10",
"11",
"10",
"00",
"10",
"00",
"01",
"11",
"01",
"01",
"00",
"01",
"00",
"00",
"11",
"11",
"00",
"01",
"11",
"01",
"00",
"10",
"11",
"00",
"11",
"10",
"01",
"00",
"00",
"00",
"10",
"11",
"10",
"11",
"10",
"10",
"00",
"00",
"10",
"11",
"01",
"00",
"10",
"11",
"01",
"01",
"01",
"11",
"10",
"01",
"10",
"01",
"10",
"00",
"10",
"01",
"00",
"00",
"01",
"10",
"01",
"11",
"11",
"10",
"11",
"10",
"11",
"11",
"10",
"01",
"11",
"00",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"01",
"11",
"11",
"10",
"01",
"11",
"01",
"10",
"00",
"00",
"00",
"10",
"00",
"01",
"10",
"11",
"10",
"11",
"00",
"11",
"01",
"11",
"10",
"11",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"01",
"00",
"01",
"00",
"00",
"11",
"00",
"01",
"11",
"00",
"10",
"10",
"10",
"11",
"11",
"00",
"00",
"10",
"10",
"11",
"01",
"01",
"01",
"01",
"11",
"11",
"00",
"11",
"00",
"01",
"01",
"10",
"01",
"11",
"00",
"11",
"10",
"01",
"01",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"11",
"11",
"11",
"01",
"10",
"01",
"00",
"10",
"00",
"11",
"00",
"00",
"10",
"00",
"01",
"01",
"00",
"10",
"11",
"10",
"01",
"11",
"01",
"10",
"11",
"11",
"01",
"10",
"11",
"10",
"01",
"00",
"01",
"00",
"01",
"10",
"10",
"01",
"11",
"01",
"11",
"11",
"10",
"00",
"00",
"11",
"10",
"00",
"11",
"00",
"00",
"11",
"10",
"00",
"11",
"11",
"01",
"01",
"01",
"10",
"01",
"11",
"00",
"01",
"10",
"11",
"10",
"10",
"11",
"11",
"00",
"00",
"11",
"10",
"01",
"01",
"11",
"11",
"10",
"10",
"00",
"00",
"10",
"01",
"10",
"00",
"01",
"11",
"00",
"11",
"11",
"11",
"10",
"11",
"11",
"11",
"01",
"10",
"00",
"01",
"10",
"10",
"01",
"10",
"01",
"10",
"00",
"01",
"11",
"01",
"00",
"10",
"11",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"10",
"00",
"10",
"11",
"11",
"01",
"01",
"11",
"10",
"10",
"10",
"11",
"11",
"11",
"00",
"10",
"11",
"01",
"11",
"11",
"01",
"10",
"01",
"10",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"11",
"00",
"00",
"01",
"10",
"11",
"11",
"00",
"00",
"00",
"00",
"11",
"00",
"11",
"11",
"10",
"10",
"10",
"11",
"11",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"01",
"10",
"00",
"11",
"00",
"00",
"00",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"10",
"11",
"10",
"01",
"01",
"00",
"00",
"11",
"01",
"10",
"11",
"10",
"10",
"01",
"11",
"00",
"11",
"10",
"00",
"10",
"01",
"00",
"01",
"10",
"10",
"11",
"01",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"11",
"00",
"01",
"00",
"11",
"10",
"00",
"00",
"10",
"00",
"00",
"01",
"00",
"00",
"01",
"00",
"00",
"11",
"10",
"01",
"11",
"10",
"11",
"00",
"00",
"10",
"10",
"10",
"00",
"01",
"10",
"10",
"10",
"11",
"01",
"11",
"10",
"00",
"10",
"01",
"00",
"11",
"00",
"10",
"01",
"11",
"00",
"00",
"00",
"01",
"01",
"10",
"11",
"01",
"01",
"10",
"01",
"11",
"10",
"10",
"01",
"01",
"00",
"11",
"11",
"00",
"00",
"11",
"01",
"10",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"11",
"11",
"01",
"00",
"10",
"01",
"00",
"01",
"11",
"00",
"11",
"00",
"11",
"00",
"00",
"00",
"11",
"01",
"00",
"01",
"00",
"10",
"11",
"11",
"10",
"10",
"11",
"10",
"00",
"00",
"11",
"10",
"00",
"01",
"01",
"00",
"01",
"01",
"01",
"00",
"11",
"10",
"01",
"10",
"00",
"11",
"00",
"00",
"11",
"11",
"00",
"10",
"11",
"11",
"01",
"10",
"01",
"11",
"01",
"01",
"11",
"01",
"00",
"00",
"11",
"11",
"01",
"11",
"01",
"00",
"10",
"01",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"01",
"01",
"00",
"11",
"01",
"11",
"01",
"01",
"11",
"00",
"00",
"00",
"10",
"10",
"01",
"00",
"01",
"10",
"11",
"11",
"00",
"11",
"11",
"01",
"11",
"10",
"10",
"00",
"11",
"00",
"11",
"01",
"00",
"11",
"01",
"01",
"10",
"00",
"10",
"01",
"11",
"11",
"00",
"10",
"01",
"00",
"10",
"01",
"00",
"00",
"01",
"11",
"10",
"01",
"11",
"01",
"01",
"01",
"01",
"10",
"01",
"11",
"10",
"00",
"10",
"10",
"10",
"00",
"11",
"11",
"11",
"10",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"00",
"01",
"01",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"10",
"00",
"11",
"11",
"00",
"01",
"00",
"11",
"11",
"11",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"01",
"01",
"11",
"01",
"10",
"01",
"01",
"01",
"01",
"10",
"00",
"10",
"01",
"10",
"01",
"00",
"00",
"10",
"10",
"01",
"01",
"00",
"01",
"01",
"00",
"01",
"00",
"11",
"11",
"01",
"10",
"01",
"10",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"10",
"10",
"11",
"00",
"01",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"00",
"11",
"01",
"01",
"11",
"00",
"10",
"11",
"00",
"00",
"10",
"00",
"00",
"11",
"01",
"00",
"00",
"01",
"01",
"00",
"11",
"11",
"00",
"00",
"01",
"00",
"01",
"10",
"00",
"10",
"01",
"00",
"11",
"10",
"00",
"10",
"00",
"01",
"10",
"11",
"01",
"00",
"00",
"10",
"01",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"01",
"00",
"10",
"00",
"01",
"10",
"11",
"11",
"00",
"00",
"01",
"11",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"01",
"00",
"11",
"10",
"01",
"11",
"11",
"01",
"11",
"01",
"01",
"11",
"11",
"10",
"10",
"10",
"00",
"00",
"10",
"00",
"11",
"11",
"10",
"01",
"00",
"10",
"01",
"00",
"11",
"01",
"01",
"11",
"10",
"00",
"11",
"01",
"01",
"01",
"10",
"11",
"10",
"00",
"11",
"01",
"11",
"10",
"00",
"10",
"01",
"10",
"10",
"11",
"11",
"01",
"10",
"00",
"00",
"11",
"00",
"11",
"10",
"11",
"01",
"00",
"10",
"00",
"11",
"11",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"10",
"01",
"01",
"10",
"11",
"10",
"11",
"11",
"01",
"10",
"10",
"11",
"10",
"00",
"00",
"10",
"00",
"11",
"10",
"01",
"11",
"10",
"00",
"00",
"00",
"00",
"10",
"01",
"10",
"01",
"01",
"11",
"00",
"01",
"00",
"00",
"00",
"11",
"11",
"00",
"10",
"00",
"10",
"00",
"10",
"10",
"11",
"00",
"01",
"10",
"00",
"10",
"01",
"11",
"10",
"01",
"10",
"01",
"10",
"01",
"11",
"10",
"11",
"00",
"11",
"00",
"11",
"10",
"00",
"01",
"10",
"00",
"00",
"10",
"10",
"01",
"01",
"00",
"00",
"01",
"01",
"11",
"11",
"01",
"00",
"01",
"00",
"00",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"10",
"01",
"10",
"10",
"01",
"11",
"10",
"10",
"01",
"10",
"00",
"01",
"11",
"00",
"11",
"00",
"01",
"10",
"11",
"01",
"00",
"11",
"00",
"10",
"00",
"01",
"10",
"00",
"11",
"01",
"10",
"11",
"00",
"01",
"00",
"11",
"11",
"01",
"11",
"00",
"10",
"11",
"10",
"11",
"01",
"11",
"11",
"11",
"10",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"01",
"10",
"01",
"10",
"01",
"00",
"10",
"10",
"01",
"10",
"00",
"10",
"01",
"10",
"01",
"01",
"00",
"10",
"01",
"10",
"10",
"01",
"00",
"00",
"00",
"11",
"10",
"11",
"10",
"01",
"00",
"00",
"01",
"11",
"00",
"11",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"01",
"01",
"11",
"11",
"00",
"01",
"10",
"00",
"11",
"11",
"00",
"10",
"11",
"00",
"10",
"10",
"00",
"11",
"10",
"11",
"10",
"10",
"11",
"00",
"00",
"10",
"10",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"10",
"00",
"11",
"01",
"00",
"00",
"01",
"10",
"11",
"11",
"10",
"11",
"00",
"01",
"01",
"11",
"10",
"00",
"01",
"10",
"00",
"11",
"01",
"01",
"10",
"11",
"11",
"10",
"11",
"00",
"10",
"10",
"01",
"01",
"11",
"01",
"10",
"00",
"01",
"10",
"11",
"11",
"00",
"11",
"01",
"11",
"10",
"10",
"10",
"11",
"01",
"11",
"00",
"00",
"00",
"00",
"01",
"00",
"10",
"11",
"01",
"00",
"10",
"11",
"01",
"11",
"00",
"00",
"10",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"01",
"01",
"10",
"10",
"00",
"00",
"10",
"01",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"00",
"11",
"01",
"10",
"11",
"00",
"10",
"00",
"10",
"01",
"00",
"11",
"11",
"00",
"10",
"10",
"00",
"00",
"10",
"00",
"11",
"10",
"01",
"01",
"00",
"10",
"00",
"01",
"01",
"01",
"10",
"00",
"11",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"00",
"01",
"01",
"01",
"10",
"00",
"01",
"11",
"11",
"10",
"10",
"11",
"10",
"11",
"11",
"10",
"11",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"11",
"11",
"01",
"11",
"00",
"01",
"01",
"11",
"01",
"01",
"00",
"00",
"00",
"00",
"01",
"10",
"01",
"00",
"10",
"00",
"11",
"10",
"01",
"11",
"00",
"01",
"00",
"11",
"00",
"00",
"10",
"11",
"00",
"10",
"11",
"11",
"00",
"01",
"11",
"01",
"10",
"00",
"10",
"00",
"01",
"11",
"11",
"00",
"10",
"10",
"01",
"11",
"00",
"01",
"11",
"00",
"11",
"01",
"10",
"11",
"11",
"00",
"10",
"01",
"00",
"10",
"00",
"01",
"01",
"11",
"11",
"00",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"10",
"00",
"10",
"10",
"11",
"11",
"01",
"00",
"10",
"11",
"00",
"10",
"01",
"01",
"11",
"10",
"10",
"11",
"00",
"11",
"01",
"10",
"01",
"10",
"11",
"10",
"10",
"11",
"00",
"11",
"00",
"00",
"01",
"11",
"11",
"10",
"01",
"10",
"01",
"11",
"11",
"11",
"01",
"00",
"00",
"01",
"01",
"10",
"01",
"01",
"10",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"01",
"10",
"00",
"00",
"01",
"01",
"00",
"01",
"10",
"11",
"00",
"11",
"01",
"00",
"10",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"10",
"10",
"00",
"01",
"11",
"10",
"10",
"10",
"10",
"10",
"01",
"00",
"00",
"00",
"10",
"00",
"11",
"10",
"10",
"10",
"00",
"11",
"01",
"01",
"00",
"01",
"01",
"10",
"00",
"11",
"10",
"00",
"01",
"11",
"11",
"10",
"01",
"11",
"10",
"10",
"00",
"10",
"00",
"01",
"11",
"00",
"10",
"00",
"01",
"01",
"10",
"00",
"01",
"10",
"10",
"11",
"00",
"00",
"11",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"00",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"01",
"01",
"00",
"01",
"11",
"11",
"10",
"10",
"00",
"10",
"00",
"01",
"00",
"10",
"11",
"01",
"01",
"01",
"11",
"01",
"01",
"10",
"00",
"01",
"11",
"01",
"10",
"10",
"11",
"11",
"11",
"10",
"10",
"10",
"01",
"00",
"01",
"10",
"11",
"01",
"10",
"00",
"10",
"10",
"11",
"00",
"00",
"10",
"00",
"01",
"01",
"11",
"10",
"10",
"00",
"00",
"00",
"11",
"10",
"10",
"11",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"11",
"10",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"10",
"00",
"00",
"11",
"01",
"01",
"11",
"01",
"00",
"11",
"00",
"01",
"10",
"00",
"01",
"10",
"01",
"10",
"00",
"00",
"11",
"11",
"11",
"11",
"10",
"00",
"00",
"00",
"10",
"11",
"10",
"10",
"00",
"01",
"11",
"01",
"01",
"01",
"11",
"00",
"00",
"01",
"10",
"11",
"11",
"01",
"10",
"01",
"01",
"00",
"00",
"01",
"10",
"10",
"01",
"01",
"11",
"00",
"10",
"10",
"10",
"00",
"01",
"11",
"10",
"11",
"10",
"00",
"00",
"01",
"00",
"11",
"10",
"11",
"01",
"11",
"01",
"10",
"10",
"10",
"01",
"01",
"10",
"11",
"00",
"00",
"11",
"00",
"10",
"10",
"10",
"01",
"01",
"11",
"01",
"10",
"11",
"00",
"10",
"11",
"10",
"01",
"11",
"10",
"10",
"10",
"10",
"01",
"00",
"11",
"01",
"11",
"00",
"00",
"11",
"00",
"00",
"10",
"10",
"00",
"11",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"10",
"01",
"10",
"11",
"10",
"01",
"11",
"00",
"00",
"11",
"01",
"01",
"11",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"11",
"01",
"00",
"01",
"01",
"10",
"00",
"00",
"10",
"10",
"10",
"01",
"11",
"01",
"01",
"01",
"01",
"11",
"10",
"11",
"10",
"11",
"00",
"11",
"01",
"01",
"11",
"00",
"00",
"01",
"10",
"11",
"11",
"11",
"10",
"00",
"01",
"10",
"11",
"00",
"11",
"11",
"00",
"11",
"00",
"01",
"10",
"10",
"10",
"10",
"10",
"00",
"11",
"01",
"10",
"01",
"01",
"10",
"00",
"00",
"11",
"10",
"01",
"01",
"10",
"10",
"00",
"11",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"11",
"00",
"11",
"10",
"00",
"11",
"10",
"01",
"11",
"00",
"11",
"11",
"10",
"00",
"01",
"01",
"01",
"00",
"11",
"11",
"00",
"00",
"00",
"00",
"11",
"11",
"01",
"10",
"00",
"00",
"01",
"10",
"00",
"10",
"11",
"01",
"01",
"00",
"10",
"11",
"01",
"10",
"11",
"11",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"11",
"00",
"11",
"01",
"11",
"10",
"10",
"11",
"01",
"00",
"10",
"00",
"11",
"10",
"11",
"10",
"10",
"10",
"01",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"01",
"00",
"00",
"10",
"10",
"11",
"11",
"01",
"10",
"11",
"00",
"01",
"01",
"11",
"00",
"01",
"10",
"10",
"00",
"10",
"01",
"10",
"10",
"01",
"00",
"10",
"11",
"10",
"11",
"00",
"01",
"11",
"10",
"11",
"10",
"00",
"11",
"11",
"11",
"00",
"01",
"11",
"00",
"01",
"10",
"01",
"01",
"01",
"10",
"10",
"00",
"00",
"11",
"00",
"01",
"00",
"10",
"00",
"11",
"11",
"10",
"01",
"00",
"11",
"01",
"00",
"01",
"10",
"10",
"00",
"01",
"10",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"10",
"00",
"10",
"11",
"10",
"11",
"10",
"00",
"00",
"01",
"01",
"10",
"01",
"11",
"11",
"00",
"10",
"10",
"01",
"01",
"00",
"01",
"01",
"11",
"01",
"11",
"11",
"00",
"01",
"01",
"00",
"11",
"10",
"01",
"10",
"01",
"00",
"10",
"10",
"11",
"11",
"00",
"00",
"00",
"01",
"00",
"01",
"10",
"00",
"10",
"10",
"10",
"11",
"10",
"00",
"01",
"11",
"01",
"01",
"10",
"00",
"10",
"10",
"00",
"10",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"00",
"11",
"10",
"10",
"01",
"10",
"00",
"01",
"10",
"11",
"10",
"00",
"00",
"00",
"10",
"10",
"10",
"11",
"10",
"10",
"01",
"11",
"00",
"01",
"01",
"01",
"00",
"01",
"10",
"10",
"11",
"00",
"11",
"00",
"01",
"00",
"00",
"01",
"01",
"00",
"11",
"10",
"00",
"11",
"11",
"01",
"00",
"00",
"01",
"10",
"01",
"01",
"00",
"00",
"10",
"10",
"10",
"11",
"00",
"11",
"01",
"11",
"11",
"11",
"00",
"00",
"01",
"10",
"11",
"11",
"10",
"10",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"00",
"10",
"10",
"01",
"10",
"10",
"01",
"01",
"01",
"11",
"11",
"00",
"01",
"10",
"10",
"01",
"01",
"11",
"10",
"00",
"01",
"11",
"10",
"10",
"00",
"01",
"10",
"00",
"00",
"01",
"10",
"11",
"00",
"10",
"10",
"00",
"10",
"11",
"10",
"00",
"00",
"11",
"01",
"11",
"01",
"00",
"00",
"10",
"01",
"11",
"01",
"00",
"11",
"10",
"11",
"00",
"00",
"11",
"11",
"11",
"01",
"10",
"00",
"00",
"01",
"01",
"10",
"01",
"00",
"11",
"11",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"00",
"01",
"10",
"11",
"00",
"10",
"01",
"10",
"11",
"10",
"00",
"00",
"11",
"00",
"01",
"11",
"10",
"00",
"10",
"10",
"11",
"11",
"00",
"10",
"01",
"10",
"00",
"10",
"00",
"00",
"10",
"11",
"00",
"00",
"01",
"01",
"00",
"00",
"00",
"11",
"11",
"00",
"10",
"00",
"00",
"11",
"01",
"00",
"10",
"11",
"10",
"00",
"01",
"01",
"01",
"10",
"01",
"01",
"00",
"01",
"00",
"10",
"11",
"10",
"01",
"11",
"01",
"10",
"11",
"00",
"11",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"10",
"10",
"10",
"11",
"11",
"00",
"10",
"01",
"11",
"10",
"01",
"10",
"01",
"00",
"11",
"01",
"00",
"11",
"01",
"01",
"00",
"10",
"10",
"11",
"11",
"01",
"01",
"11",
"01",
"11",
"00",
"00",
"01",
"01",
"00",
"00",
"11",
"10",
"11",
"10",
"11",
"01",
"11",
"01",
"10",
"10",
"10",
"01",
"01",
"00",
"10",
"11",
"10",
"01",
"11",
"11",
"01",
"01",
"11",
"10",
"01",
"11",
"01",
"01",
"10",
"10",
"10",
"01",
"11",
"11",
"01",
"00",
"00",
"10",
"10",
"10",
"01",
"11",
"10",
"00",
"11",
"10",
"11",
"10",
"00",
"00",
"00",
"11",
"01",
"01",
"10",
"10",
"00",
"01",
"10",
"11",
"11",
"01",
"10",
"11",
"10",
"00",
"00",
"01",
"01",
"10",
"01",
"11",
"11",
"11",
"00",
"00",
"10",
"11",
"11",
"10",
"11",
"11",
"11",
"00",
"10",
"00",
"11",
"00",
"01",
"00",
"10",
"10",
"11",
"10",
"10",
"01",
"00",
"10",
"00",
"10",
"11",
"10",
"00",
"00",
"11",
"01",
"01",
"01",
"11",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"01",
"01",
"00",
"01",
"10",
"01",
"10",
"10",
"11",
"10",
"11",
"00",
"10",
"11",
"10",
"11",
"10",
"01",
"10",
"00",
"01",
"00",
"10",
"01",
"00",
"00",
"01",
"00",
"11",
"00",
"10",
"10",
"00",
"10",
"00",
"10",
"00",
"01",
"01",
"10",
"01",
"00",
"01",
"10",
"10",
"11",
"01",
"01",
"11",
"10",
"01",
"10",
"10",
"00",
"00",
"01",
"10",
"01",
"11",
"11",
"00",
"10",
"10",
"10",
"10",
"11",
"11",
"01",
"01",
"01",
"10",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"01",
"11",
"11",
"11",
"00",
"11",
"00",
"00",
"01",
"11",
"10",
"11",
"00",
"10",
"11",
"00",
"00",
"01",
"11",
"11",
"11",
"11",
"00",
"01",
"01",
"11",
"01",
"10",
"10",
"00",
"11",
"11",
"11",
"10",
"00",
"10",
"11",
"11",
"01",
"00",
"01",
"10",
"11",
"11",
"11",
"10",
"11",
"11",
"11",
"01",
"01",
"11",
"01",
"00",
"01",
"01",
"01",
"00",
"00",
"10",
"10",
"10",
"00",
"01",
"00",
"01",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"11",
"00",
"11",
"10",
"01",
"00",
"10",
"01",
"11",
"00",
"00",
"00",
"10",
"00",
"00",
"00",
"10",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"01",
"01",
"01",
"10",
"11",
"10",
"11",
"10",
"11",
"00",
"00",
"11",
"01",
"01",
"01",
"01",
"00",
"10",
"01",
"01",
"10",
"11",
"00",
"01",
"11",
"10",
"00",
"00",
"00",
"11",
"11",
"01",
"00",
"10",
"00",
"00",
"01",
"01",
"11",
"00",
"10",
"10",
"10",
"11",
"11",
"10",
"00",
"01",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"10",
"00",
"01",
"10",
"00",
"11",
"11",
"00",
"01",
"00",
"00",
"00",
"10",
"01",
"00",
"11",
"00",
"01",
"11",
"10",
"11",
"11",
"11",
"11",
"10",
"10",
"00",
"00",
"00",
"10",
"10",
"01",
"00",
"11",
"11",
"00",
"11",
"10",
"01",
"01",
"11",
"01",
"00",
"10",
"01",
"01",
"00",
"00",
"10",
"01",
"11",
"01",
"00",
"10",
"11",
"11",
"10",
"00",
"11",
"01",
"01",
"00",
"00",
"11",
"00",
"01",
"10",
"11",
"01",
"01",
"11",
"11",
"11",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"11",
"01",
"10",
"10",
"01",
"00",
"00",
"10",
"00",
"01",
"10",
"10",
"01",
"01",
"01",
"01",
"11",
"11",
"00",
"11",
"01",
"11",
"01",
"11",
"00",
"01",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"10",
"00",
"11",
"10",
"01",
"11",
"00",
"10",
"00",
"00",
"01",
"00",
"11",
"11",
"01",
"10",
"00",
"00",
"11",
"00",
"01",
"01",
"11",
"01",
"11",
"10",
"10",
"00",
"11",
"00",
"01",
"11",
"10",
"01",
"00",
"01",
"00",
"11",
"11",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"00",
"01",
"01",
"01",
"00",
"11",
"00",
"11",
"01",
"00",
"10",
"10",
"11",
"01",
"10",
"00",
"11",
"01",
"01",
"00",
"11",
"00",
"11",
"01",
"00",
"11",
"01",
"01",
"01",
"00",
"11",
"01",
"10",
"00",
"01",
"11",
"00",
"01",
"01",
"00",
"00",
"01",
"11",
"11",
"01",
"00",
"10",
"01",
"10",
"00",
"11",
"11",
"00",
"11",
"10",
"00",
"11",
"11",
"00",
"10",
"01",
"01",
"00",
"11",
"10",
"00",
"10",
"01",
"11",
"01",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"10",
"01",
"01",
"00",
"00",
"01",
"10",
"11",
"01",
"01",
"10",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"01",
"00",
"00",
"10",
"11",
"11",
"01",
"01",
"10",
"01",
"01",
"00",
"10",
"11",
"00",
"11",
"11",
"00",
"00",
"01",
"00",
"11",
"00",
"11",
"00",
"00",
"10",
"10",
"10",
"10",
"00",
"00",
"11",
"11",
"00",
"00",
"11",
"10",
"10",
"00",
"00",
"11",
"01",
"01",
"01",
"10",
"11",
"11",
"10",
"01",
"11",
"01",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"01",
"10",
"11",
"10",
"00",
"01",
"11",
"10",
"11",
"10",
"01",
"10",
"01",
"10",
"00",
"11",
"11",
"11",
"01",
"11",
"00",
"11",
"11",
"00",
"01",
"01",
"01",
"11",
"10",
"00",
"01",
"10",
"00",
"11",
"00",
"00",
"00",
"11",
"10",
"11",
"11",
"10",
"10",
"11",
"11",
"10",
"10",
"10",
"11",
"00",
"00",
"01",
"00",
"11",
"10",
"10",
"10",
"01",
"11",
"10",
"00",
"00",
"01",
"00",
"01",
"01",
"00",
"10",
"01",
"10",
"10",
"00",
"11",
"00",
"00",
"11",
"10",
"10",
"00",
"01",
"00",
"01",
"10",
"00",
"01",
"11",
"00",
"00",
"00",
"11",
"11",
"11",
"10",
"11",
"10",
"10",
"01",
"01",
"00",
"01",
"10",
"11",
"01",
"00",
"10",
"11",
"00",
"00",
"01",
"00",
"01",
"00",
"11",
"10",
"00",
"11",
"00",
"10",
"10",
"11",
"11",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"10",
"01",
"11",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"11",
"00",
"01",
"01",
"00",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"01",
"00",
"11",
"01",
"01",
"11",
"11",
"10",
"11",
"10",
"01",
"10",
"01",
"11",
"00",
"11",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"01",
"00",
"10",
"01",
"10",
"00",
"01",
"00",
"01",
"10",
"01",
"00",
"01",
"11",
"01",
"01",
"00",
"10",
"10",
"10",
"10",
"01",
"00",
"11",
"00",
"10",
"00",
"00",
"00",
"11",
"10",
"10",
"10",
"10",
"10",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"10",
"00",
"10",
"00",
"01",
"01",
"11",
"11",
"11",
"00",
"01",
"11",
"11",
"10",
"11",
"00",
"00",
"00",
"10",
"10",
"00",
"11",
"10",
"10",
"11",
"00",
"10",
"00",
"01",
"10",
"01",
"01",
"01",
"00",
"11",
"11",
"00",
"00",
"10",
"10",
"10",
"11",
"00",
"10",
"01",
"11",
"00",
"00",
"10",
"00",
"00",
"10",
"10",
"01",
"01",
"11",
"11",
"01",
"10",
"00",
"01",
"01",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"10",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"11",
"00",
"10",
"00",
"10",
"10",
"11",
"01",
"10",
"00",
"11",
"10",
"10",
"10",
"00",
"10",
"10",
"00",
"00",
"00",
"01",
"00",
"10",
"10",
"00",
"00",
"10",
"11",
"11",
"00",
"11",
"01",
"11",
"01",
"10",
"01",
"11",
"10",
"00",
"10",
"10",
"01",
"01",
"00",
"01",
"01",
"00",
"01",
"01",
"00",
"00",
"10",
"00",
"11",
"11",
"01",
"00",
"01",
"10",
"11",
"10",
"10",
"00",
"00",
"11",
"11",
"01",
"01",
"11",
"10",
"00",
"10",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"01",
"11",
"10",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"01",
"01",
"01",
"01",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"11",
"11",
"11",
"01",
"10",
"00",
"01",
"11",
"11",
"00",
"10",
"01",
"10",
"00",
"11",
"01",
"10",
"00",
"01",
"10",
"01",
"11",
"10",
"01",
"10",
"11",
"10",
"00",
"10",
"11",
"11",
"11",
"00",
"11",
"01",
"00",
"00",
"11",
"10",
"10",
"01",
"00",
"01",
"11",
"10",
"10",
"11",
"00",
"11",
"00",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"01",
"01",
"11",
"10",
"10",
"00",
"00",
"01",
"10",
"11",
"10",
"10",
"00",
"00",
"01",
"11",
"01",
"11",
"00",
"01",
"00",
"01",
"10",
"11",
"00",
"01",
"10",
"00",
"11",
"11",
"01",
"01",
"01",
"11",
"00",
"10",
"10",
"10",
"10",
"10",
"10",
"11",
"00",
"11",
"01",
"01",
"11",
"11",
"10",
"11",
"10",
"01",
"11",
"11",
"01",
"11",
"11",
"01",
"00",
"00",
"11",
"10",
"01",
"00",
"11",
"10",
"11",
"10",
"01",
"11",
"10",
"00",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"10",
"10",
"11",
"00",
"01",
"11",
"11",
"01",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"01",
"01",
"00",
"10",
"00",
"10",
"01",
"01",
"11",
"11",
"11",
"11",
"00",
"01",
"01",
"10",
"00",
"00",
"10",
"11",
"11",
"10",
"00",
"01",
"00",
"01",
"11",
"00",
"00",
"11",
"10",
"11",
"00",
"10",
"11",
"10",
"00",
"00",
"00",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"00",
"00",
"11",
"01",
"00",
"11",
"00",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"01",
"11",
"00",
"01",
"11",
"00",
"11",
"10",
"00",
"01",
"01",
"01",
"11",
"11",
"10",
"00",
"01",
"01",
"00",
"01",
"00",
"01",
"01",
"10",
"11",
"00",
"01",
"11",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"00",
"00",
"00",
"10",
"01",
"10",
"10",
"11",
"11",
"01",
"11",
"10",
"00",
"00",
"11",
"00",
"11",
"10",
"11",
"10",
"01",
"01",
"10",
"00",
"00",
"11",
"10",
"00",
"10",
"01",
"10",
"01",
"10",
"00",
"00",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"10",
"10",
"10",
"01",
"10",
"10",
"10",
"10",
"00",
"01",
"11",
"11",
"01",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"11",
"11",
"00",
"10",
"01",
"10",
"10",
"10",
"01",
"10",
"01",
"11",
"01",
"01",
"11",
"10",
"00",
"00",
"01",
"01",
"11",
"11",
"00",
"01",
"11",
"00",
"10",
"11",
"10",
"00",
"00",
"10",
"10",
"10",
"11",
"01",
"00",
"11",
"11",
"01",
"11",
"10",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"00",
"01",
"10",
"10",
"10",
"00",
"01",
"11",
"11",
"01",
"01",
"01",
"11",
"01",
"11",
"00",
"10",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"10",
"11",
"11",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"10",
"11",
"11",
"00",
"11",
"10",
"01",
"00",
"01",
"10",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"11",
"10",
"00",
"01",
"01",
"11",
"11",
"11",
"00",
"00",
"00",
"00",
"11",
"10",
"01",
"01",
"10",
"10",
"01",
"10",
"10",
"01",
"10",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"00",
"01",
"00",
"00",
"11",
"10",
"01",
"11",
"00",
"11",
"01",
"10",
"01",
"10",
"10",
"01",
"00",
"10",
"11",
"11",
"10",
"11",
"00",
"01",
"10",
"00",
"00",
"01",
"11",
"00",
"00",
"01",
"10",
"10",
"01",
"11",
"10",
"00",
"01",
"10",
"00",
"00",
"11",
"01",
"01",
"01",
"00",
"11",
"11",
"01",
"01",
"11",
"10",
"01",
"11",
"11",
"11",
"10",
"01",
"10",
"10",
"00",
"10",
"00",
"00",
"01",
"10",
"10",
"01",
"01",
"01",
"11",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"01",
"10",
"00",
"11",
"01",
"11",
"10",
"00",
"10",
"00",
"11",
"10",
"01",
"11",
"11",
"11",
"11",
"01",
"10",
"00",
"01",
"00",
"10",
"10",
"00",
"00",
"01",
"11",
"01",
"01",
"00",
"00",
"01",
"11",
"01",
"00",
"01",
"00",
"00",
"11",
"00",
"10",
"01",
"01",
"01",
"11",
"10",
"10",
"00",
"01",
"01",
"11",
"01",
"01",
"01",
"11",
"10",
"01",
"01",
"10",
"11",
"11",
"00",
"11",
"10",
"11",
"00",
"10",
"01",
"11",
"11",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"01",
"00",
"10",
"11",
"00",
"01",
"10",
"10",
"11",
"10",
"11",
"10",
"10",
"00",
"11",
"00",
"01",
"01",
"11",
"01",
"01",
"11",
"10",
"10",
"00",
"01",
"10",
"00",
"01",
"11",
"11",
"01",
"01",
"10",
"11",
"01",
"01",
"10",
"01",
"11",
"10",
"01",
"01",
"11",
"11",
"01",
"00",
"11",
"01",
"10",
"11",
"00",
"01",
"00",
"10",
"10",
"01",
"00",
"00",
"01",
"10",
"00",
"01",
"00",
"10",
"10",
"11",
"10",
"01",
"11",
"10",
"01",
"11",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"00",
"01",
"01",
"00",
"01",
"01",
"00",
"01",
"00",
"11",
"00",
"10",
"00",
"00",
"11",
"01",
"01",
"00",
"11",
"11",
"00",
"01",
"00",
"10",
"01",
"10",
"01",
"01",
"10",
"00",
"01",
"11",
"00",
"11",
"10",
"11",
"00",
"10",
"01",
"11",
"01",
"01",
"10",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"00",
"10",
"00",
"11",
"11",
"11",
"11",
"10",
"00",
"01",
"11",
"11",
"10",
"10",
"11",
"00",
"00",
"10",
"11",
"10",
"00",
"10",
"01",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"10",
"01",
"00",
"00",
"10",
"00",
"00",
"11",
"11",
"10",
"00",
"01",
"01",
"10",
"11",
"01",
"10",
"11",
"00",
"01",
"11",
"01",
"10",
"11",
"10",
"00",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"01",
"00",
"00",
"01",
"00",
"00",
"10",
"01",
"00",
"00",
"10",
"10",
"01",
"10",
"01",
"10",
"01",
"10",
"01",
"00",
"10",
"00",
"00",
"10",
"00",
"01",
"00",
"11",
"00",
"11",
"11",
"01",
"00",
"10",
"11",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"01",
"10",
"11",
"00",
"00",
"10",
"00",
"10",
"11",
"11",
"01",
"11",
"01",
"10",
"00",
"11",
"11",
"10",
"11",
"10",
"00",
"10",
"01",
"01",
"10",
"10",
"11",
"11",
"00",
"00",
"11",
"01",
"10",
"00",
"10",
"10",
"11",
"00",
"01",
"10",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"01",
"11",
"10",
"11",
"01",
"11",
"01",
"00",
"10",
"01",
"00",
"01",
"00",
"00",
"01",
"10",
"00",
"11",
"11",
"01",
"01",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"00",
"11",
"00",
"01",
"10",
"00",
"10",
"01",
"11",
"01",
"00",
"01",
"00",
"11",
"01",
"11",
"11",
"01",
"00",
"00",
"01",
"10",
"10",
"00",
"00",
"01",
"10",
"00",
"01",
"00",
"00",
"10",
"10",
"00",
"10",
"11",
"00",
"10",
"10",
"10",
"00",
"00",
"00",
"10",
"01",
"01",
"00",
"00",
"00",
"10",
"00",
"01",
"10",
"00",
"01",
"01",
"01",
"00",
"01",
"10",
"11",
"10",
"01",
"00",
"00",
"11",
"10",
"01",
"01",
"10",
"10",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"01",
"00",
"11",
"10",
"11",
"00",
"00",
"11",
"00",
"10",
"10",
"01",
"00",
"00",
"00",
"11",
"11",
"01",
"11",
"00",
"10",
"00",
"01",
"10",
"01",
"10",
"01",
"10",
"10",
"11",
"00",
"01",
"00",
"00",
"10",
"01",
"00",
"01",
"10",
"00",
"10",
"10",
"11",
"11",
"11",
"10",
"11",
"11",
"11",
"00",
"00",
"01",
"11",
"10",
"01",
"11",
"11",
"11",
"01",
"11",
"01",
"01",
"10",
"00",
"10",
"00",
"01",
"11",
"01",
"01",
"00",
"00",
"10",
"00",
"00",
"10",
"01",
"00",
"00",
"01",
"00",
"10",
"01",
"00",
"11",
"01",
"00",
"00",
"01",
"10",
"11",
"10",
"10",
"11",
"00",
"11",
"01",
"10",
"01",
"01",
"10",
"01",
"00",
"01",
"01",
"01",
"11",
"00",
"00",
"11",
"10",
"10",
"00",
"11",
"10",
"00",
"00",
"00",
"11",
"11",
"10",
"01",
"00",
"11",
"01",
"10",
"00",
"10",
"00",
"11",
"11",
"01",
"01",
"11",
"00",
"10",
"01",
"11",
"10",
"00",
"00",
"10",
"11",
"00",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"11",
"01",
"00",
"11",
"11",
"11",
"00",
"10",
"00",
"00",
"00",
"00",
"11",
"10",
"01",
"10",
"00",
"11",
"01",
"10",
"00",
"01",
"00",
"11",
"10",
"11",
"11",
"11",
"11",
"01",
"00",
"00",
"00",
"11",
"00",
"11",
"01",
"10",
"10",
"01",
"11",
"11",
"00",
"00",
"01",
"01",
"10",
"10",
"11",
"11",
"00",
"11",
"01",
"11",
"10",
"10",
"00",
"01",
"00",
"11",
"11",
"10",
"00",
"11",
"01",
"00",
"00",
"10",
"01",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"01",
"10",
"11",
"00",
"00",
"00",
"01",
"01",
"10",
"01",
"11",
"01",
"10",
"10",
"00",
"01",
"11",
"01",
"01",
"11",
"00",
"10",
"11",
"10",
"10",
"10",
"00",
"11",
"00",
"10",
"10",
"11",
"00",
"01",
"00",
"00",
"00",
"01",
"10",
"01",
"11",
"11",
"11",
"11",
"11",
"11",
"11",
"01",
"10",
"11",
"11",
"01",
"00",
"10",
"11",
"00",
"01",
"11",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"11",
"01",
"00",
"10",
"01",
"00",
"01",
"10",
"11",
"00",
"11",
"01",
"00",
"11",
"11",
"11",
"11",
"11",
"01",
"11",
"10",
"00",
"10",
"10",
"10",
"11",
"01",
"01",
"01",
"10",
"01",
"11",
"11",
"01",
"11",
"10",
"00",
"11",
"01",
"10",
"00",
"11",
"11",
"00",
"00",
"00",
"11",
"01",
"00",
"10",
"01",
"00",
"00",
"01",
"00",
"10",
"10",
"00",
"01",
"01",
"00",
"00",
"01",
"11",
"10",
"11",
"10",
"10",
"00",
"11",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"10",
"01",
"11",
"11",
"00",
"11",
"11",
"01",
"00",
"01",
"10",
"01",
"10",
"01",
"11",
"01",
"11",
"00",
"10",
"10",
"01",
"11",
"11",
"10",
"10",
"10",
"00",
"00",
"01",
"10",
"01",
"01",
"01",
"10",
"11",
"11",
"00",
"01",
"00",
"11",
"11",
"00",
"10",
"10",
"01",
"11",
"01",
"00",
"11",
"10",
"11",
"01",
"10",
"10",
"01",
"11",
"10",
"00",
"10",
"00",
"10",
"01",
"01",
"00",
"01",
"11",
"11",
"10",
"01",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"10",
"01",
"10",
"00",
"01",
"11",
"00",
"01",
"00",
"00",
"00",
"00",
"01",
"01",
"10",
"11",
"00",
"10",
"01",
"10",
"10",
"01",
"10",
"01",
"01",
"01",
"11",
"11",
"10",
"10",
"10",
"11",
"11",
"00",
"11",
"01",
"10",
"10",
"11",
"11",
"00",
"00",
"00",
"10",
"11",
"10",
"10",
"00",
"10",
"00",
"10",
"10",
"01",
"11",
"11",
"01",
"10",
"00",
"10",
"10",
"01",
"11",
"10",
"01",
"10",
"00",
"10",
"11",
"01",
"01",
"01",
"10",
"11",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"11",
"01",
"11",
"10",
"11",
"00",
"00",
"11",
"11",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"01",
"00",
"01",
"10",
"00",
"01",
"00",
"00",
"01",
"11",
"01",
"00",
"11",
"11",
"11",
"10",
"01",
"10",
"10",
"00",
"00",
"00",
"01",
"00",
"10",
"00",
"00",
"01",
"10",
"00",
"01",
"11",
"00",
"10",
"01",
"00",
"01",
"11",
"00",
"10",
"01",
"00",
"01",
"11",
"10",
"01",
"10",
"01",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"10",
"10",
"10",
"00",
"00",
"01",
"11",
"10",
"00",
"01",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"01",
"10",
"01",
"11",
"10",
"00",
"10",
"10",
"11",
"00",
"01",
"00",
"00",
"11",
"00",
"10",
"00",
"10",
"10",
"11",
"01",
"10",
"01",
"10",
"10",
"01",
"11",
"11",
"00",
"11",
"11",
"00",
"11",
"11",
"11",
"10",
"01",
"10",
"00",
"01",
"11",
"10",
"10",
"00",
"11",
"10",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"00",
"10",
"01",
"10",
"00",
"01",
"00",
"01",
"00",
"11",
"01",
"11",
"01",
"11",
"00",
"10",
"01",
"11",
"01",
"10",
"11",
"10",
"11",
"10",
"01",
"00",
"00",
"01",
"10",
"00",
"01",
"00",
"11",
"00",
"01",
"11",
"01",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"00",
"00",
"01",
"01",
"01",
"01",
"00",
"01",
"01",
"11",
"01",
"01",
"10",
"00",
"11",
"00",
"01",
"11",
"10",
"01",
"10",
"11",
"01",
"10",
"00",
"11",
"01",
"01",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"01",
"00",
"00",
"01",
"00",
"00",
"00",
"01",
"11",
"01",
"01",
"10",
"11",
"00",
"01",
"01",
"00",
"11",
"00",
"10",
"00",
"10",
"01",
"10",
"01",
"11",
"11",
"01",
"01",
"10",
"11",
"00",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"11",
"00",
"00",
"00",
"10",
"01",
"00",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"10",
"00",
"01",
"10",
"10",
"01",
"10",
"01",
"11",
"10",
"11",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"00",
"01",
"11",
"00",
"00",
"01",
"00",
"00",
"01",
"11",
"01",
"11",
"01",
"01",
"00",
"01",
"00",
"00",
"00",
"10",
"01",
"11",
"01",
"10",
"11",
"00",
"00",
"00",
"00",
"10",
"10",
"01",
"11",
"01",
"10",
"01",
"10",
"01",
"00",
"01",
"01",
"10",
"00",
"00",
"10",
"01",
"00",
"10",
"11",
"10",
"01",
"10",
"00",
"10",
"00",
"00",
"10",
"00",
"10",
"11",
"00",
"00",
"10",
"00",
"10",
"11",
"10",
"11",
"00",
"10",
"01",
"00",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"01",
"11",
"00",
"00",
"10",
"01",
"10",
"00",
"11",
"01",
"11",
"00",
"01",
"01",
"00",
"11",
"11",
"01",
"00",
"00",
"10",
"11",
"10",
"11",
"10",
"10",
"11",
"00",
"01",
"01",
"01",
"10",
"11",
"10",
"10",
"11",
"11",
"11",
"00",
"11",
"10",
"00",
"00",
"11",
"00",
"11",
"11",
"01",
"10",
"10",
"00",
"10",
"11",
"00",
"11",
"10",
"11",
"01",
"00",
"01",
"11",
"01",
"00",
"00",
"01",
"11",
"10",
"01",
"00",
"10",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"01",
"01",
"10",
"00",
"10",
"00",
"00",
"01",
"00",
"11",
"10",
"01",
"10",
"00",
"11",
"00",
"11",
"01",
"01",
"01",
"10",
"01",
"00",
"10",
"11",
"10",
"01",
"00",
"01",
"11",
"10",
"11",
"00",
"00",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"00",
"10",
"01",
"01",
"10",
"11",
"01",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"01",
"01",
"10",
"00",
"01",
"01",
"11",
"11",
"10",
"10",
"11",
"11",
"01",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"00",
"01",
"11",
"10",
"01",
"01",
"01",
"00",
"10",
"00",
"10",
"01",
"01",
"00",
"10",
"11",
"10",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"00",
"10",
"00",
"10",
"10",
"00",
"10",
"11",
"01",
"10",
"11",
"00",
"01",
"11",
"10",
"00",
"00",
"10",
"11",
"01",
"01",
"00",
"01",
"01",
"01",
"10",
"01",
"10",
"11",
"10",
"11",
"11",
"10",
"00",
"10",
"00",
"10",
"00",
"10",
"01",
"11",
"00",
"10",
"11",
"10",
"00",
"01",
"10",
"00",
"10",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"11",
"00",
"01",
"01",
"10",
"00",
"01",
"01",
"00",
"11",
"01",
"01",
"00",
"00",
"11",
"10",
"11",
"11",
"11",
"11",
"01",
"10",
"00",
"11",
"11",
"00",
"10",
"01",
"00",
"11",
"11",
"10",
"01",
"11",
"11",
"10",
"00",
"11",
"00",
"01",
"10",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"01",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"10",
"00",
"01",
"00",
"11",
"01",
"10",
"00",
"01",
"01",
"00",
"01",
"11",
"00",
"10",
"01",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"00",
"00",
"10",
"11",
"00",
"11",
"01",
"11",
"00",
"11",
"01",
"10",
"10",
"11",
"10",
"11",
"00",
"01",
"11",
"01",
"00",
"00",
"01",
"00",
"10",
"11",
"10",
"11",
"00",
"11",
"01",
"11",
"00",
"11",
"01",
"01",
"00",
"01",
"11",
"00",
"01",
"00",
"00",
"11",
"11",
"01",
"10",
"10",
"11",
"00",
"01",
"01",
"11",
"11",
"01",
"10",
"00",
"00",
"10",
"11",
"01",
"10",
"01",
"11",
"00",
"11",
"00",
"10",
"00",
"11",
"01",
"01",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"10",
"00",
"00",
"01",
"11",
"10",
"01",
"11",
"11",
"11",
"01",
"11",
"01",
"00",
"00",
"11",
"00",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"01",
"10",
"10",
"01",
"00",
"01",
"00",
"00",
"01",
"00",
"01",
"00",
"00",
"10",
"00",
"10",
"11",
"10",
"01",
"11",
"10",
"01",
"01",
"10",
"10",
"00",
"00",
"10",
"10",
"11",
"11",
"10",
"10",
"10",
"11",
"01",
"10",
"01",
"10",
"11",
"01",
"10",
"01",
"10",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"00",
"00",
"00",
"01",
"00",
"10",
"11",
"11",
"10",
"00",
"10",
"00",
"10",
"00",
"00",
"01",
"01",
"10",
"00",
"00",
"10",
"01",
"10",
"01",
"01",
"01",
"01",
"10",
"01",
"01",
"01",
"11",
"01",
"10",
"11",
"11",
"10",
"11",
"10",
"10",
"01",
"10",
"00",
"01",
"01",
"00",
"10",
"01",
"00",
"01",
"00",
"11",
"11",
"11",
"10",
"10",
"00",
"01",
"01",
"01",
"00",
"11",
"01",
"00",
"11",
"10",
"00",
"10",
"10",
"11",
"00",
"00",
"11",
"01",
"10",
"01",
"01",
"01",
"00",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"00",
"10",
"11",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"01",
"00",
"01",
"10",
"11",
"11",
"01",
"10",
"00",
"10",
"11",
"01",
"00",
"11",
"01",
"10",
"10",
"01",
"10",
"10",
"11",
"10",
"01",
"11",
"11",
"00",
"00",
"01",
"11",
"00",
"10",
"01",
"01",
"10",
"10",
"00",
"01",
"01",
"11",
"01",
"00",
"10",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"01",
"01",
"00",
"10",
"11",
"01",
"10",
"01",
"10",
"00",
"00",
"00",
"11",
"00",
"01",
"01",
"01",
"01",
"10",
"01",
"11",
"00",
"10",
"00",
"11",
"11",
"01",
"11",
"00",
"01",
"11",
"10",
"00",
"01",
"10",
"01",
"00",
"11",
"01",
"10",
"01",
"11",
"01",
"01",
"00",
"11",
"01",
"10",
"00",
"10",
"00",
"01",
"11",
"11",
"00",
"01",
"00",
"01",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"10",
"01",
"11",
"01",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"10",
"00",
"00",
"01",
"10",
"11",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"11",
"10",
"01",
"01",
"11",
"00",
"00",
"10",
"11",
"11",
"11",
"00",
"10",
"11",
"01",
"01",
"00",
"11",
"10",
"11",
"10",
"10",
"11",
"10",
"00",
"11",
"01",
"11",
"00",
"10",
"11",
"00",
"10",
"10",
"10",
"00",
"11",
"11",
"10",
"01",
"10",
"00",
"11",
"11",
"00",
"01",
"11",
"00",
"10",
"00",
"11",
"10",
"11",
"01",
"01",
"11",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"00",
"11",
"01",
"01",
"00",
"10",
"10",
"11",
"11",
"00",
"01",
"11",
"11",
"00",
"10",
"00",
"11",
"00",
"01",
"01",
"00",
"10",
"11",
"10",
"10",
"00",
"01",
"10",
"01",
"00",
"11",
"11",
"11",
"10",
"10",
"01",
"00",
"11",
"11",
"00",
"00",
"11",
"00",
"01",
"10",
"10",
"01",
"00",
"01",
"00",
"10",
"10",
"01",
"01",
"10",
"11",
"11",
"01",
"10",
"11",
"11",
"01",
"11",
"10",
"11",
"10",
"01",
"00",
"10",
"01",
"01",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"10",
"00",
"00",
"01",
"11",
"01",
"01",
"00",
"10",
"01",
"11",
"01",
"01",
"01",
"00",
"01",
"11",
"11",
"01",
"10",
"00",
"11",
"10",
"10",
"11",
"11",
"11",
"00",
"10",
"00",
"10",
"11",
"01",
"11",
"11",
"11",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"10",
"00",
"01",
"10",
"11",
"11",
"00",
"00",
"10",
"01",
"11",
"11",
"00",
"00",
"01",
"01",
"11",
"00",
"11",
"00",
"01",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"00",
"00",
"11",
"10",
"10",
"10",
"10",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"10",
"10",
"01",
"00",
"00",
"11",
"11",
"11",
"01",
"10",
"00",
"01",
"01",
"11",
"00",
"10",
"01",
"00",
"10",
"00",
"11",
"01",
"01",
"11",
"01",
"10",
"10",
"00",
"00",
"00",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"11",
"00",
"10",
"11",
"00",
"11",
"01",
"00",
"01",
"00",
"11",
"01",
"10",
"00",
"01",
"11",
"01",
"11",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"00",
"11",
"11",
"10",
"00",
"10",
"10",
"10",
"11",
"10",
"00",
"11",
"00",
"10",
"01",
"01",
"10",
"00",
"11",
"11",
"00",
"01",
"11",
"01",
"00",
"11",
"01",
"10",
"00",
"10",
"01",
"10",
"11",
"00",
"00",
"10",
"11",
"00",
"10",
"11",
"10",
"11",
"01",
"10",
"10",
"00",
"01",
"10",
"10",
"10",
"10",
"01",
"00",
"10",
"11",
"10",
"00",
"11",
"00",
"00",
"00",
"11",
"01",
"11",
"01",
"10",
"10",
"11",
"10",
"01",
"11",
"10",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"00",
"10",
"01",
"10",
"11",
"10",
"01",
"11",
"01",
"01",
"11",
"01",
"00",
"01",
"11",
"01",
"00",
"11",
"10",
"11",
"01",
"01",
"10",
"11",
"00",
"10",
"10",
"11",
"00",
"11",
"00",
"00",
"11",
"01",
"11",
"10",
"00",
"00",
"11",
"10",
"10",
"11",
"11",
"10",
"10",
"00",
"10",
"01",
"10",
"11",
"10",
"01",
"00",
"00",
"00",
"10",
"10",
"10",
"01",
"10",
"01",
"10",
"00",
"01",
"00",
"11",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"01",
"01",
"10",
"10",
"11",
"01",
"10",
"00",
"01",
"10",
"01",
"00",
"00",
"10",
"00",
"10",
"11",
"00",
"01",
"10",
"11",
"10",
"01",
"11",
"11",
"01",
"01",
"01",
"10",
"00",
"11",
"10",
"01",
"10",
"10",
"10",
"01",
"11",
"00",
"00",
"11",
"11",
"11",
"11",
"10",
"10",
"00",
"01",
"11",
"01",
"00",
"00",
"00",
"01",
"10",
"11",
"11",
"00",
"11",
"00",
"01",
"01",
"01",
"00",
"11",
"01",
"01",
"00",
"00",
"11",
"10",
"01",
"11",
"11",
"01",
"11",
"11",
"00",
"01",
"00",
"01",
"11",
"01",
"10",
"10",
"11",
"00",
"01",
"01",
"10",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"00",
"00",
"11",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"01",
"11",
"10",
"10",
"10",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"00",
"01",
"10",
"11",
"10",
"11",
"01",
"11",
"11",
"00",
"11",
"00",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"10",
"10",
"01",
"00",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"01",
"10",
"10",
"10",
"10",
"10",
"00",
"01",
"11",
"10",
"10",
"00",
"00",
"10",
"11",
"01",
"11",
"11",
"11",
"01",
"01",
"01",
"00",
"10",
"11",
"00",
"11",
"11",
"10",
"01",
"11",
"11",
"01",
"11",
"10",
"11",
"01",
"10",
"10",
"01",
"01",
"11",
"11",
"00",
"00",
"11",
"00",
"00",
"01",
"10",
"00",
"11",
"11",
"01",
"10",
"01",
"00",
"11",
"00",
"11",
"10",
"00",
"10",
"10",
"00",
"10",
"00",
"11",
"10",
"01",
"10",
"01",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"01",
"10",
"00",
"00",
"00",
"11",
"10",
"10",
"01",
"00",
"11",
"11",
"10",
"00",
"00",
"11",
"11",
"10",
"01",
"10",
"01",
"10",
"11",
"11",
"10",
"01",
"10",
"11",
"00",
"11",
"00",
"11",
"01",
"11",
"10",
"11",
"10",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"10",
"11",
"11",
"01",
"11",
"11",
"10",
"01",
"11",
"10",
"10",
"01",
"00",
"01",
"01",
"01",
"10",
"01",
"01",
"11",
"10",
"10",
"00",
"00",
"10",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"01",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"00",
"10",
"10",
"01",
"01",
"11",
"00",
"01",
"00",
"11",
"11",
"01",
"11",
"11",
"01",
"11",
"10",
"11",
"00",
"10",
"11",
"11",
"00",
"11",
"10",
"10",
"11",
"11",
"00",
"10",
"00",
"00",
"11",
"00",
"11",
"10",
"11",
"00",
"10",
"11",
"11",
"01",
"10",
"01",
"00",
"11",
"00",
"01",
"00",
"01",
"01",
"10",
"10",
"11",
"00",
"01",
"10",
"10",
"01",
"10",
"00",
"11",
"00",
"00",
"01",
"11",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"00",
"10",
"01",
"11",
"00",
"00",
"11",
"01",
"01",
"00",
"11",
"10",
"11",
"10",
"10",
"01",
"11",
"01",
"01",
"11",
"01",
"00",
"11",
"10",
"11",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"11",
"01",
"01",
"10",
"11",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"01",
"11",
"01",
"01",
"01",
"11",
"01",
"00",
"10",
"10",
"01",
"00",
"11",
"00",
"00",
"01",
"00",
"00",
"11",
"00",
"00",
"11",
"00",
"11",
"01",
"10",
"10",
"00",
"00",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"11",
"10",
"01",
"10",
"11",
"10",
"00",
"01",
"01",
"10",
"00",
"00",
"01",
"00",
"01",
"01",
"00",
"11",
"01",
"11",
"00",
"11",
"11",
"00",
"11",
"10",
"01",
"11",
"11",
"10",
"11",
"01",
"00",
"00",
"01",
"11",
"10",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"00",
"11",
"00",
"10",
"01",
"11",
"11",
"01",
"00",
"01",
"10",
"01",
"11",
"01",
"01",
"01",
"00",
"11",
"11",
"11",
"10",
"10",
"10",
"11",
"10",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"01",
"00",
"00",
"00",
"00",
"11",
"10",
"10",
"10",
"01",
"00",
"11",
"00",
"11",
"10",
"01",
"01",
"00",
"00",
"00",
"11",
"10",
"11",
"11",
"00",
"10",
"10",
"01",
"10",
"10",
"11",
"10",
"00",
"01",
"01",
"11",
"10",
"11",
"10",
"10",
"11",
"11",
"01",
"00",
"00",
"01",
"11",
"01",
"00",
"11",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"00",
"10",
"10",
"01",
"01",
"11",
"01",
"01",
"10",
"11",
"11",
"10",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"10",
"00",
"00",
"10",
"01",
"00",
"10",
"10",
"10",
"10",
"01",
"11",
"11",
"11",
"00",
"00",
"00",
"10",
"11",
"11",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"11",
"11",
"01",
"10",
"01",
"10",
"01",
"00",
"00",
"10",
"10",
"00",
"00",
"01",
"11",
"10",
"00",
"10",
"10",
"01",
"10",
"00",
"11",
"01",
"01",
"11",
"11",
"10",
"01",
"10",
"10",
"10",
"11",
"01",
"01",
"01",
"10",
"11",
"00",
"00",
"10",
"10",
"00",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"01",
"11",
"01",
"11",
"01",
"11",
"00",
"11",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"10",
"01",
"10",
"11",
"11",
"01",
"00",
"01",
"01",
"10",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"11",
"11",
"10",
"00",
"11",
"00",
"11",
"01",
"01",
"00",
"01",
"00",
"00",
"10",
"00",
"10",
"11",
"00",
"00",
"10",
"10",
"11",
"10",
"00",
"01",
"11",
"01",
"01",
"01",
"00",
"11",
"10",
"00",
"01",
"11",
"00",
"10",
"00",
"11",
"00",
"01",
"01",
"00",
"11",
"00",
"10",
"01",
"10",
"11",
"00",
"01",
"11",
"11",
"00",
"01",
"00",
"11",
"11",
"00",
"00",
"10",
"10",
"01",
"11",
"00",
"11",
"10",
"10",
"00",
"01",
"01",
"00",
"00",
"10",
"10",
"00",
"11",
"11",
"00",
"11",
"00",
"11",
"11",
"01",
"11",
"00",
"00",
"11",
"00",
"00",
"11",
"10",
"01",
"00",
"10",
"10",
"00",
"11",
"11",
"11",
"11",
"11",
"10",
"11",
"01",
"00",
"01",
"11",
"10",
"11",
"10",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"00",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"11",
"10",
"11",
"01",
"01",
"01",
"01",
"10",
"11",
"11",
"10",
"01",
"00",
"11",
"11",
"10",
"00",
"10",
"11",
"11",
"00",
"00",
"10",
"00",
"01",
"01",
"00",
"00",
"10",
"00",
"01",
"11",
"01",
"00",
"00",
"01",
"00",
"00",
"01",
"01",
"00",
"00",
"10",
"11",
"10",
"11",
"11",
"00",
"00",
"00",
"01",
"11",
"11",
"01",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"00",
"01",
"00",
"11",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"01",
"00",
"00",
"00",
"10",
"00",
"01",
"01",
"10",
"00",
"10",
"00",
"10",
"10",
"11",
"10",
"11",
"10",
"01",
"01",
"01",
"00",
"10",
"00",
"00",
"10",
"10",
"00",
"00",
"10",
"01",
"00",
"01",
"00",
"00",
"00",
"11",
"11",
"00",
"00",
"00",
"10",
"11",
"10",
"01",
"11",
"00",
"11",
"00",
"00",
"11",
"10",
"11",
"10",
"10",
"01",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"11",
"00",
"11",
"00",
"00",
"00",
"11",
"00",
"11",
"00",
"11",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"00",
"00",
"10",
"10",
"01",
"01",
"01",
"01",
"01",
"10",
"01",
"10",
"01",
"01",
"00",
"00",
"11",
"11",
"00",
"10",
"11",
"10",
"11",
"01",
"00",
"11",
"00",
"11",
"11",
"00",
"01",
"01",
"10",
"11",
"11",
"10",
"00",
"01",
"11",
"00",
"00",
"00",
"10",
"00",
"10",
"10",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"01",
"11",
"11",
"11",
"10",
"10",
"11",
"11",
"10",
"10",
"01",
"11",
"01",
"10",
"11",
"11",
"11",
"00",
"00",
"10",
"10",
"10",
"11",
"11",
"11",
"10",
"00",
"01",
"10",
"11",
"10",
"01",
"01",
"01",
"00",
"11",
"11",
"00",
"10",
"00",
"00",
"01",
"10",
"10",
"00",
"11",
"11",
"10",
"11",
"11",
"10",
"11",
"11",
"01",
"11",
"10",
"10",
"10",
"11",
"11",
"00",
"01",
"00",
"01",
"01",
"00",
"01",
"11",
"10",
"10",
"11",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"00",
"00",
"00",
"11",
"00",
"10",
"11",
"00",
"00",
"00",
"11",
"10",
"10",
"00",
"11",
"11",
"11",
"10",
"01",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"10",
"00",
"11",
"10",
"11",
"11",
"00",
"01",
"00",
"01",
"10",
"00",
"00",
"11",
"01",
"00",
"10",
"00",
"10",
"10",
"01",
"01",
"00",
"01",
"01",
"00",
"10",
"11",
"10",
"00",
"11",
"10",
"10",
"00",
"11",
"10",
"00",
"11",
"11",
"11",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"01",
"11",
"11",
"01",
"10",
"10",
"11",
"00",
"10",
"11",
"00",
"00",
"11",
"00",
"11",
"01",
"00",
"11",
"11",
"00",
"00",
"00",
"00",
"10",
"01",
"11",
"11",
"10",
"01",
"10",
"00",
"10",
"11",
"00",
"11",
"00",
"11",
"00",
"11",
"11",
"00",
"10",
"10",
"00",
"00",
"00",
"10",
"10",
"10",
"11",
"00",
"11",
"11",
"01",
"10",
"11",
"00",
"01",
"01",
"00",
"10",
"10",
"11",
"11",
"00",
"11",
"00",
"10",
"00",
"10",
"01",
"10",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"11",
"11",
"10",
"10",
"01",
"11",
"11",
"00",
"00",
"00",
"00",
"11",
"10",
"10",
"11",
"11",
"01",
"00",
"11",
"00",
"10",
"11",
"00",
"10",
"01",
"00",
"11",
"10",
"00",
"10",
"10",
"11",
"01",
"11",
"11",
"10",
"11",
"11",
"00",
"11",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"11",
"11",
"01",
"11",
"11",
"01",
"10",
"11",
"00",
"10",
"00",
"10",
"00",
"01",
"10",
"11",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"00",
"10",
"11",
"00",
"10",
"01",
"11",
"01",
"01",
"10",
"00",
"00",
"00",
"11",
"00",
"00",
"01",
"00",
"11",
"11",
"00",
"00",
"01",
"00",
"00",
"00",
"01",
"01",
"10",
"01",
"10",
"11",
"11",
"00",
"10",
"00",
"11",
"10",
"11",
"01",
"11",
"01",
"10",
"10",
"00",
"10",
"00",
"10",
"10",
"00",
"00",
"11",
"10",
"01",
"11",
"10",
"11",
"10",
"10",
"00",
"00",
"10",
"00",
"10",
"00",
"01",
"11",
"10",
"00",
"01",
"10",
"00",
"10",
"00",
"00",
"11",
"00",
"10",
"01",
"11",
"00",
"11",
"01",
"11",
"00",
"01",
"00",
"00",
"01",
"00",
"11",
"10",
"00",
"01",
"10",
"00",
"01",
"11",
"01",
"11",
"01",
"00",
"10",
"11",
"00",
"11",
"00",
"00",
"01",
"11",
"01",
"01",
"00",
"11",
"11",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"00",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"00",
"11",
"10",
"01",
"10",
"10",
"11",
"11",
"11",
"10",
"10",
"00",
"01",
"01",
"00",
"01",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"00",
"11",
"10",
"10",
"01",
"00",
"01",
"10",
"11",
"10",
"00",
"10",
"11",
"01",
"00",
"01",
"10",
"11",
"01",
"00",
"10",
"00",
"11",
"01",
"11",
"00",
"10",
"01",
"01",
"00",
"10",
"11",
"00",
"01",
"01",
"10",
"10",
"11",
"10",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"10",
"10",
"10",
"11",
"01",
"10",
"11",
"00",
"00",
"00",
"01",
"10",
"10",
"01",
"00",
"00",
"01",
"01",
"01",
"11",
"11",
"10",
"10",
"00",
"00",
"01",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"01",
"00",
"00",
"00",
"11",
"01",
"01",
"11",
"00",
"10",
"00",
"11",
"00",
"11",
"01",
"01",
"11",
"01",
"00",
"01",
"01",
"11",
"00",
"00",
"11",
"10",
"00",
"00",
"01",
"00",
"11",
"01",
"00",
"00",
"00",
"01",
"10",
"10",
"00",
"01",
"10",
"01",
"10",
"10",
"11",
"01",
"10",
"00",
"10",
"00",
"10",
"10",
"00",
"11",
"01",
"01",
"00",
"00",
"00",
"11",
"00",
"01",
"01",
"01",
"01",
"11",
"10",
"11",
"01",
"00",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"01",
"00",
"00",
"10",
"01",
"01",
"00",
"10",
"00",
"00",
"10",
"01",
"10",
"11",
"00",
"00",
"01",
"10",
"01",
"00",
"00",
"01",
"11",
"00",
"00",
"10",
"11",
"11",
"00",
"01",
"11",
"10",
"10",
"01",
"01",
"00",
"00",
"01",
"10",
"11",
"01",
"10",
"01",
"10",
"10",
"10",
"01",
"01",
"00",
"01",
"01",
"00",
"01",
"01",
"00",
"00",
"10",
"00",
"11",
"01",
"10",
"00",
"01",
"11",
"00",
"10",
"10",
"00",
"00",
"11",
"11",
"01",
"11",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"11",
"10",
"11",
"10",
"10",
"11",
"00",
"01",
"11",
"11",
"00",
"00",
"00",
"00",
"01",
"00",
"11",
"01",
"00",
"11",
"01",
"00",
"00",
"10",
"11",
"00",
"00",
"01",
"00",
"01",
"10",
"10",
"00",
"00",
"11",
"00",
"11",
"10",
"11",
"10",
"01",
"10",
"01",
"00",
"11",
"10",
"00",
"01",
"10",
"01",
"11",
"10",
"11",
"11",
"00",
"11",
"01",
"11",
"00",
"01",
"01",
"01",
"11",
"01",
"00",
"11",
"00",
"00",
"01",
"11",
"00",
"11",
"00",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"10",
"00",
"11",
"00",
"10",
"11",
"11",
"00",
"10",
"10",
"11",
"00",
"00",
"01",
"01",
"10",
"11",
"00",
"00",
"00",
"11",
"01",
"11",
"10",
"10",
"11",
"00",
"10",
"01",
"10",
"10",
"11",
"01",
"10",
"10",
"11",
"00",
"01",
"00",
"00",
"01",
"11",
"01",
"00",
"00",
"10",
"11",
"10",
"11",
"10",
"00",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"01",
"11",
"00",
"10",
"00",
"11",
"00",
"01",
"01",
"01",
"11",
"11",
"00",
"01",
"10",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"00",
"11",
"01",
"10",
"10",
"00",
"10",
"00",
"10",
"10",
"00",
"01",
"01",
"00",
"01",
"10",
"10",
"10",
"11",
"00",
"00",
"11",
"01",
"10",
"00",
"11",
"10",
"11",
"01",
"01",
"01",
"11",
"10",
"01",
"01",
"00",
"01",
"00",
"01",
"00",
"00",
"01",
"00",
"10",
"01",
"00",
"11",
"11",
"00",
"11",
"10",
"10",
"00",
"10",
"01",
"00",
"11",
"01",
"10",
"10",
"01",
"00",
"11",
"11",
"00",
"11",
"10",
"00",
"00",
"00",
"11",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"10",
"01",
"11",
"01",
"00",
"10",
"11",
"00",
"00",
"00",
"10",
"00",
"01",
"01",
"11",
"10",
"00",
"00",
"10",
"00",
"11",
"01",
"10",
"01",
"11",
"01",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"00",
"00",
"11",
"10",
"10",
"10",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"10",
"00",
"01",
"01",
"00",
"00",
"01",
"11",
"11",
"11",
"01",
"11",
"10",
"01",
"01",
"11",
"11",
"00",
"11",
"01",
"01",
"10",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"00",
"10",
"01",
"10",
"11",
"11",
"11",
"10",
"00",
"11",
"01",
"01",
"00",
"00",
"10",
"01",
"00",
"00",
"01",
"10",
"11",
"11",
"01",
"11",
"11",
"00",
"11",
"01",
"00",
"00",
"00",
"11",
"11",
"10",
"10",
"00",
"11",
"11",
"11",
"01",
"00",
"10",
"01",
"01",
"10",
"10",
"11",
"00",
"11",
"00",
"11",
"10",
"10",
"01",
"11",
"01",
"00",
"01",
"10",
"11",
"00",
"10",
"00",
"10",
"10",
"00",
"11",
"00",
"10",
"01",
"10",
"00",
"11",
"01",
"00",
"00",
"11",
"10",
"10",
"00",
"10",
"10",
"11",
"01",
"10",
"00",
"00",
"11",
"11",
"01",
"10",
"00",
"11",
"00",
"11",
"11",
"00",
"01",
"10",
"01",
"00",
"01",
"11",
"00",
"10",
"00",
"11",
"10",
"10",
"00",
"01",
"00",
"11",
"01",
"01",
"00",
"11",
"01",
"11",
"11",
"01",
"00",
"10",
"11",
"10",
"01",
"11",
"11",
"10",
"01",
"10",
"10",
"01",
"11",
"01",
"00",
"11",
"10",
"00",
"10",
"10",
"10",
"00",
"01",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"10",
"10",
"10",
"00",
"01",
"00",
"11",
"00",
"01",
"11",
"10",
"11",
"11",
"01",
"00",
"11",
"11",
"01",
"10",
"00",
"10",
"10",
"00",
"11",
"11",
"10",
"11",
"10",
"11",
"11",
"01",
"01",
"00",
"11",
"01",
"11",
"00",
"00",
"10",
"00",
"11",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"10",
"00",
"00",
"00",
"11",
"00",
"00",
"00",
"11",
"10",
"00",
"11",
"11",
"10",
"10",
"01",
"10",
"00",
"10",
"11",
"10",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"01",
"00",
"00",
"01",
"10",
"10",
"10",
"01",
"01",
"01",
"01",
"01",
"01",
"01",
"11",
"10",
"00",
"11",
"00",
"11",
"11",
"10",
"01",
"01",
"10",
"10",
"10",
"10",
"11",
"10",
"01",
"00",
"11",
"01",
"10",
"00",
"11",
"00",
"10",
"10",
"00",
"10",
"00",
"00",
"11",
"01",
"01",
"11",
"00",
"10",
"11",
"10",
"01",
"10",
"10",
"01",
"11",
"11",
"01",
"10",
"11",
"11",
"10",
"00",
"11",
"10",
"10",
"10",
"10",
"11",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"10",
"10",
"10",
"10",
"00",
"00",
"11",
"10",
"01",
"01",
"00",
"10",
"11",
"00",
"10",
"10",
"11",
"01",
"00",
"01",
"11",
"00",
"11",
"10",
"10",
"00",
"10",
"10",
"10",
"10",
"11",
"11",
"00",
"01",
"10",
"00",
"00",
"11",
"11",
"10",
"01",
"01",
"01",
"00",
"01",
"10",
"11",
"00",
"11",
"00",
"01",
"10",
"10",
"10",
"10",
"11",
"11",
"10",
"11",
"11",
"01",
"00",
"11",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"01",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"01",
"10",
"01",
"11",
"01",
"01",
"01",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"10",
"01",
"00",
"00",
"01",
"00",
"11",
"00",
"01",
"10",
"00",
"00",
"01",
"01",
"00",
"11",
"01",
"10",
"01",
"11",
"10",
"10",
"00",
"11",
"00",
"10",
"11",
"01",
"11",
"00",
"11",
"11",
"10",
"00",
"01",
"01",
"01",
"00",
"10",
"01",
"01",
"11",
"00",
"00",
"11",
"11",
"11",
"10",
"00",
"01",
"11",
"00",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"01",
"00",
"10",
"11",
"00",
"10",
"01",
"00",
"00",
"00",
"01",
"11",
"11",
"10",
"00",
"10",
"01",
"11",
"01",
"10",
"01",
"10",
"00",
"10",
"11",
"10",
"11",
"00",
"01",
"00",
"01",
"11",
"11",
"00",
"10",
"11",
"01",
"00",
"01",
"00",
"01",
"10",
"10",
"00",
"10",
"01",
"10",
"01",
"01",
"11",
"01",
"01",
"11",
"01",
"11",
"10",
"11",
"10",
"01",
"00",
"01",
"00",
"10",
"10",
"01",
"11",
"10",
"10",
"10",
"00",
"10",
"01",
"10",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"00",
"10",
"00",
"01",
"01",
"00",
"00",
"01",
"00",
"11",
"00",
"10",
"01",
"00",
"11",
"11",
"01",
"10",
"11",
"11",
"00",
"10",
"01",
"00",
"00",
"11",
"10",
"01",
"10",
"10",
"10",
"11",
"01",
"00",
"00",
"00",
"11",
"10",
"01",
"10",
"11",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"01",
"11",
"10",
"11",
"11",
"11",
"00",
"00",
"01",
"01",
"00",
"01",
"11",
"00",
"11",
"10",
"11",
"11",
"10",
"00",
"01",
"11",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"10",
"01",
"10",
"01",
"01",
"11",
"00",
"10",
"00",
"10",
"00",
"01",
"11",
"01",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"01",
"00",
"00",
"00",
"10",
"00",
"10",
"11",
"00",
"11",
"10",
"11",
"01",
"01",
"00",
"00",
"11",
"10",
"01",
"10",
"01",
"10",
"00",
"01",
"11",
"01",
"11",
"00",
"00",
"01",
"10",
"11",
"11",
"10",
"10",
"11",
"01",
"11",
"10",
"00",
"00",
"10",
"10",
"11",
"10",
"11",
"01",
"11",
"00",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"00",
"10",
"00",
"01",
"01",
"01",
"10",
"11",
"01",
"01",
"10",
"00",
"00",
"11",
"00",
"01",
"01",
"00",
"00",
"10",
"10",
"11",
"01",
"10",
"00",
"00",
"11",
"11",
"10",
"10",
"10",
"10",
"10",
"11",
"00",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"10",
"11",
"11",
"00",
"01",
"11",
"01",
"10",
"00",
"00",
"11",
"11",
"00",
"10",
"10",
"10",
"11",
"00",
"11",
"01",
"11",
"11",
"01",
"10",
"01",
"10",
"11",
"00",
"00",
"00",
"11",
"00",
"01",
"01",
"11",
"10",
"01",
"00",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"01",
"00",
"11",
"11",
"00",
"00",
"10",
"10",
"01",
"01",
"01",
"10",
"00",
"10",
"11",
"00",
"00",
"00",
"11",
"01",
"10",
"01",
"11",
"00",
"11",
"01",
"01",
"10",
"01",
"00",
"00",
"00",
"10",
"11",
"00",
"00",
"01",
"11",
"00",
"10",
"11",
"11",
"00",
"10",
"10",
"11",
"10",
"10",
"10",
"01",
"11",
"01",
"01",
"11",
"11",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"01",
"01",
"01",
"00",
"01",
"10",
"11",
"00",
"01",
"01",
"11",
"00",
"00",
"00",
"10",
"10",
"10",
"11",
"11",
"01",
"01",
"00",
"00",
"00",
"00",
"11",
"10",
"00",
"01",
"00",
"00",
"10",
"10",
"10",
"11",
"10",
"01",
"01",
"10",
"11",
"10",
"00",
"10",
"01",
"11",
"01",
"00",
"01",
"01",
"00",
"00",
"10",
"00",
"01",
"10",
"10",
"00",
"01",
"01",
"10",
"00",
"11",
"01",
"11",
"00",
"01",
"11",
"01",
"10",
"10",
"00",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"11",
"10",
"00",
"01",
"10",
"11",
"11",
"01",
"10",
"11",
"01",
"11",
"01",
"00",
"10",
"10",
"00",
"11",
"00",
"11",
"10",
"01",
"10",
"10",
"00",
"11",
"00",
"10",
"10",
"01",
"00",
"10",
"00",
"01",
"00",
"10",
"10",
"00",
"00",
"10",
"10",
"11",
"11",
"01",
"00",
"10",
"11",
"11",
"10",
"01",
"11",
"10",
"10",
"10",
"10",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"00",
"11",
"01",
"11",
"11",
"01",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"11",
"10",
"10",
"11",
"11",
"10",
"00",
"10",
"11",
"10",
"00",
"11",
"01",
"11",
"10",
"00",
"11",
"11",
"11",
"11",
"11",
"00",
"11",
"01",
"01",
"11",
"00",
"10",
"01",
"00",
"11",
"10",
"00",
"01",
"01",
"11",
"00",
"11",
"00",
"10",
"10",
"01",
"00",
"01",
"10",
"00",
"10",
"00",
"01",
"01",
"01",
"00",
"01",
"01",
"00",
"10",
"10",
"00",
"00",
"10",
"00",
"11",
"11",
"00",
"10",
"10",
"11",
"10",
"01",
"10",
"01",
"11",
"10",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"01",
"00",
"01",
"11",
"01",
"00",
"00",
"00",
"00",
"01",
"00",
"00",
"10",
"01",
"01",
"01",
"00",
"10",
"10",
"11",
"10",
"11",
"10",
"00",
"00",
"11",
"11",
"11",
"10",
"00",
"11",
"00",
"01",
"01",
"10",
"10",
"00",
"01",
"10",
"00",
"10",
"01",
"00",
"01",
"10",
"11",
"10",
"10",
"01",
"10",
"01",
"11",
"11",
"01",
"10",
"11",
"10",
"11",
"01",
"10",
"00",
"01",
"10",
"01",
"10",
"00",
"01",
"11",
"01",
"11",
"11",
"01",
"10",
"10",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"00",
"01",
"11",
"10",
"10",
"01",
"00",
"00",
"01",
"11",
"11",
"00",
"10",
"01",
"11",
"00",
"11",
"00",
"10",
"01",
"10",
"10",
"10",
"11",
"11",
"10",
"01",
"00",
"11",
"00",
"10",
"00",
"11",
"01",
"11",
"01",
"01",
"00",
"01",
"11",
"10",
"00",
"00",
"00",
"11",
"00",
"00",
"11",
"01",
"11",
"10",
"00",
"01",
"00",
"01",
"10",
"01",
"10",
"11",
"00",
"10",
"10",
"00",
"11",
"11",
"00",
"10",
"11",
"01",
"10",
"10",
"00",
"11",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"10",
"01",
"11",
"11",
"00",
"00",
"11",
"10",
"01",
"00",
"10",
"10",
"00",
"11",
"01",
"01",
"01",
"01",
"00",
"10",
"00",
"11",
"11",
"00",
"00",
"01",
"01",
"00",
"10",
"11",
"10",
"10",
"10",
"11",
"00",
"00",
"00",
"01",
"01",
"11",
"00",
"11",
"10",
"10",
"00",
"10",
"00",
"01",
"10",
"10",
"00",
"00",
"11",
"00",
"10",
"11",
"00",
"01",
"11",
"10",
"00",
"00",
"01",
"11",
"01",
"01",
"10",
"11",
"10",
"11",
"00",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"11",
"11",
"01",
"10",
"11",
"00",
"00",
"10",
"10",
"00",
"11",
"10",
"00",
"00",
"00",
"11",
"10",
"10",
"00",
"11",
"00",
"10",
"00",
"10",
"01",
"00",
"01",
"01",
"00",
"01",
"10",
"01",
"00",
"11",
"11",
"00",
"10",
"10",
"00",
"11",
"10",
"11",
"00",
"00",
"11",
"11",
"01",
"11",
"11",
"10",
"10",
"10",
"10",
"11",
"10",
"00",
"01",
"01",
"00",
"11",
"01",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"11",
"11",
"11",
"11",
"00",
"01",
"10",
"01",
"10",
"01",
"10",
"01",
"00",
"00",
"00",
"11",
"10",
"01",
"00",
"11",
"00",
"01",
"10",
"10",
"11",
"00",
"11",
"00",
"11",
"11",
"01",
"00",
"00",
"10",
"00",
"10",
"11",
"10",
"00",
"10",
"01",
"10",
"01",
"01",
"10",
"01",
"00",
"10",
"01",
"00",
"11",
"11",
"11",
"00",
"01",
"10",
"01",
"11",
"11",
"00",
"10",
"00",
"00",
"10",
"11",
"11",
"10",
"11",
"10",
"01",
"01",
"10",
"01",
"11",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"11",
"10",
"00",
"01",
"00",
"11",
"01",
"01",
"00",
"00",
"10",
"01",
"10",
"01",
"00",
"00",
"10",
"00",
"11",
"11",
"01",
"11",
"11",
"00",
"00",
"01",
"10",
"01",
"11",
"10",
"10",
"10",
"11",
"11",
"10",
"00",
"01",
"11",
"10",
"11",
"00",
"00",
"00",
"10",
"11",
"01",
"01",
"10",
"11",
"00",
"10",
"10",
"00",
"11",
"11",
"00",
"10",
"10",
"11",
"10",
"10",
"10",
"01",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"10",
"11",
"10",
"11",
"01",
"01",
"00",
"00",
"01",
"10",
"10",
"01",
"00",
"00",
"11",
"11",
"00",
"01",
"01",
"10",
"10",
"10",
"00",
"00",
"00",
"11",
"10",
"10",
"11",
"10",
"10",
"01",
"11",
"10",
"11",
"11",
"10",
"11",
"10",
"01",
"00",
"00",
"01",
"11",
"00",
"01",
"11",
"01",
"10",
"01",
"01",
"00",
"10",
"00",
"11",
"10",
"00",
"11",
"11",
"00",
"00",
"00",
"10",
"00",
"01",
"11",
"01",
"10",
"10",
"11",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"00",
"01",
"10",
"11",
"11",
"11",
"01",
"00",
"00",
"10",
"00",
"11",
"00",
"00",
"00",
"11",
"00",
"01",
"01",
"11",
"00",
"00",
"00",
"00",
"10",
"00",
"00",
"10",
"11",
"01",
"10",
"00",
"11",
"01",
"11",
"10",
"00",
"00",
"01",
"01",
"11",
"10",
"01",
"01",
"01",
"10",
"11",
"01",
"11",
"01",
"11",
"10",
"00",
"11",
"01",
"11",
"11",
"00",
"00",
"11",
"10",
"01",
"01",
"00",
"00",
"11",
"00",
"11",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"10",
"11",
"01",
"10",
"11",
"10",
"01",
"01",
"00",
"11",
"00",
"01",
"01",
"01",
"00",
"01",
"01",
"01",
"11",
"00",
"01",
"10",
"11",
"11",
"10",
"01",
"10",
"01",
"11",
"10",
"00",
"00",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"01",
"00",
"01",
"11",
"10",
"10",
"01",
"00",
"01",
"00",
"11",
"00",
"10",
"10",
"00",
"01",
"01",
"00",
"10",
"11",
"01",
"10",
"00",
"10",
"10",
"10",
"00",
"11",
"11",
"11",
"10",
"01",
"11",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"10",
"11",
"10",
"01",
"10",
"11",
"01",
"11",
"11",
"01",
"01",
"10",
"11",
"11",
"01",
"01",
"10",
"01",
"11",
"11",
"00",
"11",
"01",
"11",
"10",
"00",
"10",
"00",
"11",
"01",
"10",
"00",
"10",
"00",
"00",
"11",
"00",
"11",
"00",
"10",
"11",
"11",
"01",
"10",
"00",
"01",
"10",
"10",
"10",
"10",
"10",
"00",
"11",
"10",
"11",
"11",
"00",
"00",
"11",
"01",
"00",
"01",
"00",
"00",
"00",
"11",
"01",
"11",
"10",
"10",
"10",
"10",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"01",
"10",
"10",
"11",
"10",
"00",
"00",
"01",
"00",
"10",
"11",
"00",
"01",
"00",
"00",
"00",
"01",
"10",
"01",
"00",
"11",
"11",
"01",
"11",
"01",
"01",
"00",
"10",
"11",
"10",
"10",
"10",
"01",
"10",
"10",
"01",
"01",
"01",
"01",
"11",
"01",
"00",
"00",
"11",
"00",
"11",
"10",
"01",
"00",
"01",
"11",
"10",
"10",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"01",
"10",
"10",
"10",
"01",
"01",
"00",
"00",
"11",
"10",
"11",
"11",
"11",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"00",
"10",
"11",
"01",
"00",
"01",
"00",
"11",
"00",
"10",
"11",
"01",
"10",
"10",
"01",
"01",
"10",
"01",
"11",
"00",
"11",
"01",
"11",
"00",
"11",
"10",
"10",
"00",
"00",
"11",
"01",
"11",
"00",
"01",
"10",
"01",
"00",
"01",
"01",
"10",
"11",
"00",
"01",
"10",
"11",
"01",
"10",
"10",
"11",
"00",
"11",
"10",
"00",
"01",
"01",
"00",
"10",
"01",
"01",
"10",
"10",
"10",
"11",
"10",
"11",
"11",
"00",
"01",
"01",
"11",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"11",
"01",
"01",
"01",
"01",
"11",
"10",
"00",
"10",
"11",
"00",
"10",
"01",
"11",
"00",
"00",
"11",
"10",
"10",
"11",
"00",
"01",
"10",
"01",
"11",
"00",
"11",
"00",
"00",
"10",
"11",
"10",
"10",
"00",
"10",
"00",
"00",
"11",
"01",
"10",
"10",
"10",
"11",
"10",
"01",
"01",
"01",
"11",
"11",
"10",
"00",
"10",
"00",
"11",
"10",
"11",
"11",
"00",
"00",
"11",
"11",
"01",
"10",
"11",
"11",
"10",
"01",
"11",
"01",
"11",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"10",
"10",
"10",
"10",
"00",
"10",
"00",
"00",
"00",
"01",
"11",
"11",
"00",
"00",
"00",
"10",
"11",
"11",
"10",
"11",
"01",
"00",
"11",
"01",
"11",
"00",
"11",
"10",
"10",
"11",
"00",
"10",
"00",
"11",
"11",
"11",
"01",
"01",
"11",
"00",
"00",
"11",
"10",
"11",
"11",
"01",
"10",
"01",
"10",
"01",
"00",
"01",
"00",
"00",
"11",
"10",
"10",
"01",
"01",
"10",
"00",
"01",
"01",
"00",
"01",
"11",
"10",
"10",
"10",
"01",
"01",
"10",
"00",
"11",
"10",
"10",
"01",
"01",
"00",
"11",
"01",
"10",
"11",
"01",
"11",
"01",
"00",
"01",
"11",
"00",
"01",
"00",
"00",
"10",
"00",
"00",
"11",
"00",
"11",
"11",
"01",
"11",
"10",
"10",
"10",
"10",
"10",
"11",
"11",
"01",
"01",
"10",
"10",
"10",
"00",
"10",
"11",
"00",
"10",
"11",
"01",
"10",
"00",
"10",
"11",
"01",
"10",
"11",
"01",
"10",
"01",
"10",
"01",
"01",
"10",
"00",
"10",
"00",
"11",
"00",
"10",
"11",
"10",
"00",
"01",
"00",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"00",
"10",
"00",
"10",
"11",
"10",
"11",
"00",
"00",
"10",
"10",
"01",
"11",
"10",
"01",
"01",
"01",
"01",
"01",
"00",
"11",
"01",
"01",
"00",
"00",
"00",
"01",
"00",
"11",
"11",
"01",
"00",
"10",
"01",
"01",
"01",
"01",
"11",
"11",
"11",
"00",
"00",
"01",
"01",
"10",
"11",
"00",
"10",
"01",
"11",
"00",
"00",
"10",
"10",
"01",
"01",
"00",
"10",
"01",
"01",
"00",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"00",
"11",
"01",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"01",
"00",
"10",
"00",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"01",
"00",
"01",
"11",
"11",
"11",
"00",
"00",
"00",
"01",
"11",
"10",
"00",
"00",
"10",
"10",
"10",
"11",
"01",
"01",
"10",
"10",
"01",
"10",
"00",
"11",
"00",
"01",
"10",
"11",
"01",
"10",
"01",
"01",
"00",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"01",
"01",
"11",
"00",
"10",
"01",
"01",
"11",
"00",
"10",
"10",
"00",
"11",
"11",
"10",
"01",
"10",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"00",
"10",
"01",
"00",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"10",
"00",
"00",
"11",
"00",
"11",
"10",
"01",
"11",
"00",
"00",
"11",
"00",
"00",
"00",
"00",
"11",
"00",
"10",
"01",
"11",
"11",
"01",
"11",
"01",
"01",
"11",
"10",
"10",
"11",
"11",
"00",
"10",
"10",
"01",
"01",
"10",
"11",
"11",
"01",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"00",
"10",
"00",
"00",
"01",
"10",
"01",
"01",
"10",
"01",
"00",
"01",
"00",
"11",
"01",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"11",
"00",
"00",
"00",
"11",
"01",
"10",
"10",
"00",
"01",
"10",
"10",
"00",
"01",
"01",
"00",
"11",
"11",
"10",
"01",
"10",
"10",
"01",
"01",
"01",
"00",
"01",
"11",
"00",
"10",
"00",
"11",
"11",
"11",
"11",
"00",
"00",
"11",
"10",
"11",
"00",
"11",
"10",
"00",
"11",
"10",
"01",
"00",
"11",
"00",
"11",
"10",
"10",
"10",
"00",
"11",
"00",
"00",
"00",
"00",
"01",
"11",
"11",
"01",
"00",
"11",
"00",
"10",
"10",
"01",
"01",
"10",
"00",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"00",
"11",
"10",
"01",
"01",
"11",
"10",
"00",
"11",
"00",
"10",
"11",
"11",
"01",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"00",
"01",
"10",
"10",
"01",
"10",
"01",
"10",
"10",
"01",
"11",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"11",
"00",
"11",
"01",
"00",
"11",
"10",
"11",
"01",
"11",
"10",
"01",
"11",
"10",
"00",
"01",
"01",
"01",
"01",
"11",
"10",
"11",
"00",
"11",
"11",
"11",
"00",
"01",
"00",
"11",
"01",
"11",
"01",
"11",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"01",
"01",
"10",
"10",
"10",
"10",
"11",
"10",
"10",
"11",
"11",
"11",
"01",
"01",
"00",
"10",
"11",
"11",
"00",
"10",
"10",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"00",
"01",
"00",
"10",
"01",
"01",
"11",
"10",
"00",
"01",
"01",
"11",
"00",
"11",
"00",
"01",
"01",
"10",
"00",
"10",
"00",
"11",
"11",
"01",
"10",
"00",
"00",
"11",
"00",
"01",
"01",
"11",
"00",
"10",
"11",
"01",
"11",
"00",
"01",
"10",
"11",
"01",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"01",
"01",
"01",
"11",
"00",
"01",
"01",
"10",
"11",
"10",
"11",
"11",
"10",
"11",
"11",
"10",
"00",
"11",
"10",
"01",
"00",
"01",
"10",
"00",
"11",
"11",
"01",
"01",
"01",
"11",
"00",
"10",
"10",
"10",
"10",
"11",
"00",
"11",
"00",
"01",
"00",
"00",
"11",
"00",
"10",
"10",
"10",
"11",
"10",
"00",
"11",
"11",
"00",
"10",
"00",
"10",
"00",
"11",
"10",
"11",
"11",
"01",
"11",
"00",
"01",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"11",
"10",
"01",
"11",
"01",
"11",
"00",
"01",
"11",
"01",
"01",
"01",
"10",
"00",
"10",
"10",
"00",
"01",
"01",
"11",
"11",
"11",
"10",
"01",
"10",
"10",
"11",
"00",
"01",
"10",
"10",
"11",
"10",
"10",
"11",
"11",
"01",
"10",
"11",
"01",
"10",
"11",
"01",
"00",
"11",
"01",
"10",
"01",
"00",
"00",
"01",
"01",
"10",
"11",
"01",
"00",
"11",
"10",
"10",
"00",
"10",
"10",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"01",
"11",
"10",
"00",
"11",
"01",
"11",
"01",
"11",
"00",
"11",
"01",
"10",
"01",
"10",
"11",
"00",
"01",
"11",
"11",
"10",
"01",
"11",
"01",
"01",
"01",
"11",
"10",
"11",
"10",
"10",
"11",
"00",
"11",
"01",
"11",
"01",
"01",
"10",
"10",
"11",
"00",
"10",
"10",
"11",
"10",
"01",
"00",
"00",
"11",
"01",
"01",
"00",
"01",
"01",
"00",
"01",
"10",
"10",
"11",
"00",
"11",
"00",
"10",
"10",
"11",
"11",
"11",
"10",
"11",
"10",
"11",
"00",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"01",
"10",
"10",
"00",
"11",
"10",
"00",
"01",
"10",
"00",
"11",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"00",
"00",
"11",
"00",
"00",
"01",
"11",
"11",
"01",
"11",
"01",
"01",
"01",
"10",
"10",
"00",
"11",
"01",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"11",
"10",
"10",
"11",
"01",
"10",
"01",
"11",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"10",
"01",
"11",
"00",
"00",
"10",
"01",
"01",
"01",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"01",
"00",
"01",
"00",
"11",
"11",
"10",
"10",
"10",
"10",
"10",
"00",
"00",
"00",
"10",
"01",
"01",
"00",
"01",
"01",
"11",
"11",
"00",
"10",
"01",
"01",
"10",
"11",
"10",
"00",
"01",
"10",
"11",
"01",
"10",
"10",
"10",
"00",
"11",
"01",
"01",
"11",
"10",
"00",
"01",
"01",
"11",
"00",
"01",
"11",
"01",
"10",
"01",
"11",
"01",
"00",
"00",
"01",
"10",
"11",
"11",
"10",
"01",
"10",
"11",
"11",
"00",
"11",
"11",
"11",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"10",
"10",
"01",
"10",
"11",
"01",
"11",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"00",
"01",
"01",
"10",
"00",
"11",
"00",
"11",
"00",
"00",
"01",
"01",
"00",
"00",
"10",
"00",
"01",
"00",
"11",
"10",
"00",
"01",
"11",
"10",
"00",
"01",
"11",
"01",
"01",
"10",
"11",
"01",
"00",
"10",
"00",
"00",
"10",
"00",
"11",
"10",
"01",
"10",
"11",
"10",
"00",
"10",
"01",
"10",
"01",
"10",
"10",
"11",
"11",
"11",
"10",
"01",
"11",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"10",
"10",
"00",
"10",
"01",
"01",
"11",
"00",
"00",
"00",
"11",
"10",
"10",
"01",
"11",
"01",
"00",
"01",
"10",
"10",
"11",
"11",
"11",
"00",
"01",
"11",
"11",
"00",
"10",
"00",
"01",
"01",
"01",
"10",
"11",
"11",
"01",
"01",
"11",
"11",
"01",
"00",
"10",
"00",
"01",
"10",
"11",
"11",
"11",
"10",
"10",
"00",
"10",
"00",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"10",
"01",
"00",
"00",
"01",
"01",
"11",
"11",
"11",
"00",
"01",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"11",
"10",
"11",
"00",
"11",
"01",
"00",
"11",
"11",
"00",
"10",
"01",
"01",
"11",
"10",
"01",
"00",
"00",
"11",
"00",
"10",
"11",
"10",
"01",
"10",
"11",
"10",
"11",
"01",
"01",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"11",
"01",
"10",
"11",
"00",
"01",
"00",
"10",
"11",
"00",
"00",
"00",
"10",
"10",
"00",
"10",
"00",
"10",
"00",
"00",
"00",
"10",
"01",
"11",
"01",
"11",
"11",
"10",
"10",
"01",
"00",
"01",
"01",
"11",
"01",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"10",
"11",
"00",
"00",
"00",
"01",
"11",
"01",
"10",
"11",
"00",
"00",
"10",
"00",
"01",
"00",
"00",
"00",
"01",
"00",
"00",
"11",
"11",
"10",
"00",
"01",
"01",
"01",
"01",
"00",
"01",
"01",
"11",
"01",
"11",
"10",
"01",
"00",
"11",
"00",
"11",
"01",
"00",
"01",
"10",
"10",
"00",
"11",
"10",
"11",
"00",
"01",
"10",
"11",
"11",
"00",
"01",
"10",
"11",
"11",
"11",
"01",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"10",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"11",
"00",
"11",
"10",
"11",
"10",
"00",
"10",
"00",
"00",
"00",
"11",
"00",
"11",
"10",
"01",
"01",
"11",
"01",
"11",
"11",
"10",
"01",
"00",
"10",
"10",
"11",
"11",
"01",
"01",
"01",
"01",
"00",
"01",
"01",
"00",
"10",
"11",
"11",
"11",
"01",
"01",
"00",
"10",
"01",
"11",
"11",
"00",
"01",
"10",
"10",
"10",
"10",
"01",
"01",
"10",
"10",
"11",
"00",
"11",
"10",
"11",
"00",
"00",
"01",
"01",
"10",
"01",
"00",
"10",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"10",
"10",
"10",
"11",
"11",
"10",
"01",
"01",
"00",
"11",
"10",
"11",
"01",
"00",
"00",
"10",
"01",
"11",
"11",
"00",
"00",
"00",
"01",
"10",
"11",
"11",
"00",
"11",
"11",
"01",
"11",
"11",
"01",
"11",
"00",
"00",
"11",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"10",
"00",
"11",
"11",
"01",
"00",
"00",
"10",
"01",
"11",
"00",
"10",
"11",
"11",
"11",
"00",
"01",
"10",
"11",
"00",
"00",
"10",
"00",
"11",
"11",
"00",
"11",
"11",
"10",
"00",
"11",
"01",
"00",
"01",
"11",
"10",
"00",
"11",
"11",
"01",
"10",
"11",
"00",
"10",
"10",
"00",
"01",
"10",
"11",
"11",
"10",
"00",
"10",
"00",
"10",
"10",
"00",
"10",
"11",
"00",
"10",
"11",
"10",
"01",
"01",
"00",
"10",
"00",
"10",
"01",
"00",
"11",
"00",
"10",
"00",
"10",
"11",
"00",
"00",
"10",
"10",
"00",
"01",
"11",
"01",
"10",
"11",
"11",
"01",
"11",
"01",
"01",
"00",
"11",
"10",
"00",
"00",
"11",
"01",
"01",
"01",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"00",
"01",
"01",
"11",
"01",
"10",
"00",
"10",
"01",
"11",
"00",
"11",
"00",
"00",
"11",
"10",
"00",
"01",
"00",
"00",
"00",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"10",
"10",
"01",
"00",
"11",
"01",
"00",
"11",
"11",
"10",
"10",
"11",
"11",
"01",
"11",
"10",
"10",
"10",
"11",
"00",
"00",
"00",
"00",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"00",
"10",
"10",
"10",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"10",
"00",
"00",
"01",
"01",
"10",
"11",
"10",
"11",
"10",
"11",
"11",
"01",
"00",
"11",
"01",
"11",
"01",
"00",
"01",
"10",
"01",
"10",
"10",
"01",
"00",
"01",
"10",
"11",
"11",
"10",
"10",
"00",
"11",
"10",
"01",
"01",
"00",
"10",
"11",
"10",
"00",
"01",
"01",
"10",
"00",
"10",
"11",
"11",
"00",
"10",
"10",
"11",
"01",
"01",
"01",
"11",
"10",
"01",
"01",
"01",
"10",
"01",
"01",
"11",
"11",
"01",
"10",
"11",
"10",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"01",
"11",
"01",
"10",
"10",
"00",
"01",
"11",
"00",
"00",
"01",
"00",
"11",
"01",
"00",
"00",
"01",
"00",
"11",
"01",
"10",
"01",
"11",
"10",
"01",
"11",
"10",
"00",
"11",
"11",
"00",
"10",
"10",
"00",
"00",
"01",
"10",
"00",
"10",
"11",
"11",
"00",
"10",
"11",
"11",
"11",
"11",
"01",
"10",
"10",
"11",
"00",
"01",
"00",
"10",
"10",
"00",
"00",
"10",
"01",
"01",
"00",
"01",
"01",
"11",
"00",
"10",
"00",
"10",
"11",
"10",
"10",
"01",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"00",
"00",
"01",
"10",
"01",
"11",
"10",
"10",
"10",
"01",
"00",
"10",
"11",
"10",
"01",
"10",
"10",
"10",
"11",
"11",
"00",
"10",
"01",
"01",
"11",
"00",
"11",
"00",
"00",
"11",
"10",
"00",
"01",
"11",
"11",
"10",
"01",
"01",
"10",
"10",
"11",
"00",
"11",
"10",
"00",
"11",
"11",
"00",
"11",
"10",
"00",
"10",
"00",
"01",
"11",
"11",
"00",
"01",
"01",
"11",
"01",
"01",
"00",
"00",
"01",
"10",
"11",
"00",
"10",
"10",
"11",
"00",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"11",
"01",
"11",
"11",
"00",
"10",
"00",
"01",
"01",
"11",
"00",
"01",
"01",
"10",
"11",
"01",
"00",
"11",
"10",
"11",
"01",
"11",
"01",
"11",
"01",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"00",
"10",
"01",
"01",
"10",
"01",
"01",
"00",
"00",
"11",
"00",
"11",
"00",
"11",
"00",
"00",
"11",
"11",
"01",
"01",
"00",
"01",
"10",
"10",
"01",
"11",
"10",
"00",
"01",
"01",
"00",
"01",
"00",
"11",
"10",
"01",
"11",
"00",
"01",
"01",
"10",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"10",
"11",
"01",
"10",
"10",
"01",
"01",
"10",
"01",
"10",
"01",
"11",
"00",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"01",
"11",
"10",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"01",
"01",
"11",
"11",
"10",
"01",
"11",
"00",
"01",
"11",
"11",
"00",
"01",
"00",
"00",
"10",
"00",
"01",
"01",
"11",
"11",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"11",
"11",
"00",
"00",
"11",
"10",
"11",
"10",
"01",
"01",
"11",
"11",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"01",
"11",
"10",
"11",
"01",
"01",
"10",
"10",
"11",
"01",
"10",
"10",
"00",
"00",
"11",
"01",
"11",
"00",
"11",
"00",
"11",
"01",
"01",
"11",
"10",
"11",
"10",
"01",
"11",
"01",
"10",
"10",
"10",
"10",
"11",
"00",
"00",
"01",
"11",
"10",
"01",
"01",
"11",
"10",
"10",
"01",
"10",
"11",
"01",
"00",
"11",
"01",
"10",
"10",
"01",
"10",
"11",
"01",
"00",
"01",
"10",
"00",
"10",
"00",
"10",
"00",
"11",
"11",
"00",
"11",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"01",
"00",
"11",
"00",
"00",
"00",
"01",
"01",
"10",
"01",
"11",
"10",
"00",
"00",
"00",
"10",
"01",
"11",
"00",
"11",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"01",
"11",
"10",
"10",
"01",
"00",
"10",
"01",
"10",
"11",
"01",
"01",
"10",
"00",
"01",
"11",
"01",
"10",
"10",
"01",
"10",
"00",
"00",
"11",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"01",
"10",
"11",
"10",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"11",
"00",
"11",
"00",
"10",
"10",
"01",
"00",
"01",
"01",
"11",
"01",
"00",
"11",
"11",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"10",
"00",
"00",
"11",
"01",
"01",
"00",
"01",
"10",
"10",
"11",
"11",
"00",
"00",
"10",
"01",
"11",
"10",
"10",
"01",
"11",
"00",
"01",
"11",
"11",
"00",
"01",
"00",
"01",
"00",
"00",
"01",
"10",
"01",
"00",
"10",
"01",
"01",
"10",
"01",
"10",
"01",
"00",
"10",
"01",
"01",
"01",
"00",
"00",
"01",
"11",
"11",
"10",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"10",
"11",
"01",
"11",
"01",
"00",
"01",
"10",
"00",
"11",
"00",
"00",
"11",
"00",
"11",
"11",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"00",
"01",
"10",
"01",
"11",
"00",
"00",
"11",
"10",
"10",
"11",
"11",
"10",
"00",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"10",
"00",
"00",
"10",
"01",
"00",
"10",
"00",
"01",
"11",
"10",
"00",
"01",
"01",
"11",
"00",
"01",
"00",
"11",
"01",
"11",
"11",
"00",
"01",
"10",
"01",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"10",
"11",
"10",
"01",
"00",
"11",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"01",
"10",
"10",
"01",
"01",
"11",
"01",
"00",
"10",
"01",
"01",
"00",
"11",
"11",
"01",
"01",
"00",
"01",
"01",
"01",
"10",
"00",
"00",
"01",
"01",
"01",
"11",
"00",
"10",
"11",
"01",
"10",
"00",
"00",
"10",
"01",
"10",
"11",
"10",
"01",
"00",
"11",
"11",
"01",
"00",
"10",
"10",
"11",
"11",
"01",
"10",
"10",
"00",
"01",
"01",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"00",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"00",
"00",
"01",
"01",
"10",
"01",
"00",
"00",
"00",
"01",
"10",
"00",
"11",
"00",
"01",
"11",
"10",
"00",
"10",
"00",
"00",
"11",
"10",
"10",
"11",
"11",
"01",
"00",
"11",
"00",
"00",
"01",
"10",
"01",
"01",
"00",
"00",
"01",
"01",
"00",
"01",
"11",
"00",
"11",
"11",
"11",
"11",
"01",
"11",
"11",
"11",
"00",
"10",
"01",
"01",
"11",
"01",
"00",
"10",
"00",
"11",
"11",
"01",
"10",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"10",
"01",
"00",
"00",
"11",
"01",
"11",
"01",
"00",
"00",
"01",
"00",
"11",
"01",
"10",
"01",
"01",
"00",
"01",
"01",
"11",
"10",
"10",
"01",
"00",
"10",
"11",
"00",
"00",
"10",
"01",
"00",
"00",
"10",
"11",
"10",
"11",
"10",
"10",
"10",
"00",
"01",
"01",
"00",
"10",
"10",
"00",
"11",
"10",
"00",
"00",
"01",
"00",
"00",
"01",
"11",
"11",
"01",
"01",
"01",
"01",
"00",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"01",
"11",
"10",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"01",
"01",
"11",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"10",
"00",
"11",
"00",
"01",
"10",
"00",
"00",
"00",
"01",
"01",
"11",
"10",
"11",
"10",
"01",
"00",
"00",
"01",
"11",
"10",
"00",
"01",
"01",
"01",
"10",
"11",
"00",
"11",
"10",
"00",
"00",
"10",
"01",
"00",
"11",
"00",
"00",
"00",
"00",
"01",
"10",
"11",
"11",
"00",
"10",
"01",
"01",
"01",
"01",
"00",
"01",
"00",
"11",
"11",
"11",
"10",
"11",
"01",
"01",
"01",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"00",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"10",
"11",
"01",
"00",
"01",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"11",
"01",
"11",
"00",
"01",
"10",
"10",
"10",
"01",
"11",
"10",
"10",
"01",
"00",
"10",
"10",
"00",
"00",
"01",
"11",
"01",
"11",
"11",
"10",
"10",
"10",
"00",
"11",
"10",
"01",
"11",
"01",
"11",
"11",
"00",
"00",
"10",
"01",
"11",
"10",
"11",
"11",
"01",
"00",
"00",
"01",
"10",
"11",
"00",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"10",
"10",
"00",
"00",
"01",
"01",
"00",
"11",
"11",
"01",
"10",
"00",
"11",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"10",
"00",
"01",
"11",
"10",
"11",
"00",
"11",
"11",
"01",
"11",
"01",
"01",
"01",
"10",
"00",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"00",
"00",
"00",
"11",
"01",
"00",
"01",
"11",
"01",
"00",
"10",
"00",
"10",
"10",
"11",
"01",
"11",
"10",
"00",
"10",
"10",
"01",
"10",
"01",
"11",
"11",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"01",
"11",
"00",
"10",
"11",
"00",
"00",
"11",
"10",
"10",
"00",
"00",
"10",
"00",
"00",
"00",
"01",
"00",
"11",
"11",
"10",
"01",
"01",
"01",
"01",
"11",
"01",
"11",
"00",
"11",
"01",
"01",
"10",
"00",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"01",
"11",
"10",
"01",
"11",
"10",
"11",
"10",
"01",
"00",
"01",
"00",
"00",
"10",
"10",
"11",
"10",
"01",
"10",
"00",
"11",
"11",
"00",
"00",
"01",
"01",
"10",
"11",
"10",
"00",
"01",
"11",
"01",
"00",
"10",
"01",
"10",
"01",
"11",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"11",
"11",
"00",
"00",
"11",
"00",
"11",
"00",
"10",
"01",
"10",
"00",
"11",
"01",
"11",
"01",
"01",
"11",
"01",
"00",
"11",
"11",
"01",
"11",
"10",
"10",
"10",
"10",
"00",
"00",
"01",
"00",
"01",
"00",
"10",
"11",
"01",
"10",
"00",
"01",
"01",
"10",
"11",
"11",
"01",
"01",
"10",
"01",
"11",
"10",
"11",
"11",
"01",
"10",
"00",
"10",
"01",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"01",
"00",
"00",
"00",
"10",
"10",
"00",
"11",
"10",
"00",
"01",
"01",
"00",
"10",
"10",
"11",
"01",
"00",
"10",
"10",
"01",
"11",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"00",
"10",
"01",
"00",
"11",
"11",
"10",
"00",
"11",
"00",
"11",
"10",
"11",
"10",
"11",
"10",
"10",
"00",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"01",
"01",
"11",
"11",
"00",
"00",
"00",
"00",
"10",
"10",
"01",
"11",
"11",
"11",
"11",
"01",
"01",
"01",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"01",
"00",
"10",
"00",
"11",
"10",
"10",
"11",
"10",
"11",
"10",
"00",
"10",
"01",
"11",
"11",
"01",
"00",
"10",
"01",
"00",
"10",
"11",
"01",
"00",
"11",
"11",
"01",
"00",
"00",
"01",
"01",
"00",
"11",
"01",
"01",
"11",
"00",
"01",
"00",
"11",
"00",
"11",
"10",
"10",
"01",
"00",
"10",
"11",
"10",
"11",
"10",
"10",
"00",
"10",
"10",
"01",
"11",
"01",
"10",
"11",
"10",
"01",
"00",
"10",
"00",
"11",
"01",
"01",
"01",
"11",
"00",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"00",
"10",
"01",
"11",
"00",
"01",
"01",
"00",
"01",
"11",
"11",
"00",
"00",
"01",
"01",
"00",
"10",
"01",
"01",
"10",
"00",
"01",
"01",
"11",
"00",
"01",
"11",
"00",
"11",
"10",
"01",
"11",
"11",
"10",
"10",
"00",
"10",
"00",
"10",
"01",
"01",
"10",
"11",
"00",
"11",
"01",
"10",
"00",
"00",
"11",
"00",
"00",
"11",
"00",
"10",
"11",
"00",
"11",
"01",
"11",
"00",
"01",
"11",
"00",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"00",
"11",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"00",
"00",
"10",
"01",
"11",
"01",
"01",
"00",
"00",
"11",
"10",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"00",
"00",
"01",
"01",
"11",
"10",
"01",
"11",
"10",
"10",
"11",
"00",
"11",
"01",
"10",
"11",
"10",
"11",
"10",
"10",
"10",
"10",
"11",
"11",
"00",
"11",
"01",
"11",
"11",
"11",
"00",
"01",
"00",
"01",
"01",
"11",
"00",
"10",
"01",
"11",
"11",
"11",
"10",
"01",
"01",
"00",
"00",
"00",
"11",
"11",
"00",
"10",
"01",
"01",
"01",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"00",
"10",
"01",
"01",
"01",
"00",
"00",
"01",
"10",
"10",
"01",
"11",
"10",
"01",
"10",
"01",
"00",
"10",
"01",
"00",
"10",
"10",
"11",
"11",
"11",
"10",
"00",
"01",
"10",
"10",
"00",
"00",
"10",
"11",
"00",
"11",
"01",
"01",
"11",
"01",
"10",
"00",
"00",
"10",
"01",
"11",
"01",
"11",
"00",
"10",
"00",
"10",
"11",
"11",
"00",
"01",
"11",
"11",
"00",
"00",
"01",
"01",
"00",
"10",
"00",
"11",
"11",
"11",
"10",
"01",
"01",
"11",
"11",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"01",
"01",
"11",
"11",
"00",
"00",
"11",
"10",
"01",
"11",
"11",
"11",
"01",
"10",
"01",
"00",
"00",
"10",
"01",
"01",
"11",
"00",
"10",
"11",
"10",
"01",
"00",
"01",
"01",
"11",
"00",
"00",
"00",
"00",
"10",
"01",
"11",
"11",
"11",
"10",
"11",
"11",
"01",
"00",
"01",
"10",
"10",
"10",
"10",
"11",
"01",
"11",
"00",
"11",
"11",
"10",
"01",
"01",
"10",
"00",
"00",
"11",
"10",
"10",
"01",
"11",
"01",
"10",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"01",
"01",
"00",
"01",
"00",
"00",
"10",
"00",
"11",
"11",
"10",
"00",
"11",
"01",
"11",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"01",
"11",
"00",
"01",
"01",
"00",
"01",
"00",
"01",
"10",
"10",
"00",
"00",
"00",
"01",
"10",
"01",
"10",
"11",
"01",
"10",
"11",
"00",
"10",
"10",
"00",
"00",
"01",
"10",
"11",
"10",
"10",
"10",
"01",
"10",
"01",
"10",
"00",
"11",
"00",
"10",
"11",
"11",
"10",
"11",
"11",
"01",
"10",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"01",
"11",
"01",
"01",
"11",
"01",
"01",
"00",
"11",
"01",
"01",
"00",
"01",
"00",
"00",
"01",
"01",
"11",
"10",
"00",
"10",
"11",
"01",
"11",
"01",
"00",
"10",
"11",
"00",
"00",
"01",
"01",
"11",
"10",
"01",
"10",
"00",
"00",
"11",
"10",
"01",
"01",
"00",
"11",
"11",
"00",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"10",
"11",
"00",
"00",
"00",
"11",
"11",
"11",
"01",
"11",
"10",
"00",
"10",
"00",
"10",
"11",
"01",
"11",
"01",
"11",
"10",
"01",
"00",
"01",
"10",
"10",
"01",
"10",
"11",
"10",
"00",
"11",
"01",
"00",
"00",
"00",
"11",
"11",
"01",
"11",
"01",
"10",
"00",
"01",
"10",
"10",
"00",
"01",
"11",
"10",
"11",
"00",
"00",
"11",
"11",
"00",
"01",
"00",
"00",
"01",
"10",
"00",
"01",
"10",
"01",
"10",
"01",
"01",
"01",
"00",
"01",
"11",
"01",
"11",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"00",
"01",
"10",
"01",
"01",
"10",
"01",
"11",
"01",
"00",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"01",
"01",
"10",
"10",
"10",
"10",
"00",
"10",
"00",
"00",
"11",
"11",
"00",
"00",
"10",
"00",
"10",
"10",
"11",
"00",
"00",
"10",
"11",
"11",
"00",
"00",
"01",
"11",
"01",
"10",
"00",
"01",
"00",
"00",
"10",
"10",
"11",
"10",
"10",
"11",
"10",
"00",
"00",
"10",
"10",
"01",
"10",
"01",
"10",
"11",
"10",
"10",
"10",
"10",
"01",
"10",
"00",
"10",
"11",
"11",
"11",
"10",
"11",
"10",
"11",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"11",
"00",
"10",
"11",
"10",
"10",
"01",
"11",
"00",
"11",
"11",
"00",
"00",
"01",
"10",
"11",
"11",
"01",
"10",
"11",
"01",
"01",
"01",
"00",
"11",
"10",
"11",
"10",
"00",
"10",
"10",
"00",
"00",
"11",
"01",
"00",
"11",
"00",
"11",
"00",
"00",
"10",
"10",
"10",
"00",
"01",
"01",
"00",
"10",
"00",
"11",
"11",
"11",
"01",
"01",
"11",
"10",
"01",
"10",
"10",
"01",
"00",
"11",
"00",
"01",
"00",
"10",
"11",
"10",
"11",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"11",
"00",
"00",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"00",
"11",
"11",
"00",
"00",
"10",
"01",
"10",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"01",
"00",
"01",
"00",
"01",
"00",
"10",
"00",
"11",
"00",
"10",
"11",
"01",
"10",
"10",
"11",
"10",
"11",
"11",
"11",
"10",
"00",
"01",
"01",
"00",
"01",
"01",
"01",
"11",
"11",
"10",
"01",
"00",
"11",
"01",
"00",
"11",
"11",
"10",
"01",
"01",
"00",
"01",
"01",
"10",
"10",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"00",
"01",
"10",
"00",
"10",
"00",
"00",
"10",
"11",
"10",
"10",
"00",
"00",
"01",
"01",
"10",
"00",
"00",
"10",
"00",
"11",
"11",
"01",
"00",
"01",
"11",
"00",
"00",
"11",
"00",
"11",
"01",
"10",
"11",
"01",
"01",
"01",
"00",
"00",
"11",
"10",
"01",
"10",
"00",
"01",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"11",
"10",
"01",
"00",
"01",
"11",
"10",
"00",
"11",
"11",
"00",
"00",
"01",
"10",
"10",
"01",
"01",
"00",
"01",
"01",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"10",
"01",
"01",
"01",
"11",
"01",
"00",
"11",
"10",
"11",
"01",
"11",
"01",
"11",
"10",
"01",
"01",
"00",
"00",
"10",
"00",
"01",
"00",
"10",
"10",
"10",
"00",
"00",
"00",
"10",
"11",
"00",
"10",
"01",
"01",
"11",
"11",
"11",
"11",
"11",
"01",
"01",
"00",
"10",
"01",
"00",
"11",
"01",
"10",
"00",
"11",
"00",
"10",
"11",
"00",
"01",
"01",
"01",
"01",
"11",
"11",
"00",
"01",
"00",
"01",
"11",
"10",
"11",
"10",
"11",
"00",
"11",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"01",
"10",
"11",
"01",
"10",
"01",
"11",
"11",
"11",
"01",
"10",
"01",
"01",
"10",
"11",
"00",
"11",
"00",
"10",
"00",
"10",
"01",
"00",
"01",
"11",
"10",
"11",
"01",
"01",
"10",
"10",
"00",
"10",
"00",
"11",
"10",
"10",
"01",
"00",
"01",
"01",
"10",
"00",
"00",
"00",
"11",
"01",
"00",
"00",
"00",
"11",
"11",
"01",
"11",
"10",
"00",
"11",
"11",
"10",
"00",
"01",
"11",
"00",
"11",
"10",
"11",
"10",
"11",
"01",
"11",
"11",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"01",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"11",
"10",
"01",
"11",
"11",
"10",
"00",
"11",
"11",
"10",
"00",
"10",
"11",
"10",
"00",
"11",
"10",
"11",
"11",
"01",
"00",
"10",
"00",
"00",
"01",
"11",
"00",
"00",
"11",
"11",
"01",
"11",
"01",
"10",
"01",
"10",
"01",
"01",
"10",
"00",
"01",
"11",
"00",
"10",
"01",
"01",
"10",
"10",
"01",
"11",
"01",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"11",
"11",
"10",
"11",
"01",
"00",
"10",
"10",
"00",
"11",
"11",
"00",
"01",
"10",
"01",
"00",
"10",
"10",
"01",
"00",
"00",
"01",
"11",
"11",
"00",
"01",
"00",
"10",
"00",
"11",
"10",
"11",
"10",
"01",
"01",
"01",
"11",
"01",
"11",
"01",
"00",
"11",
"00",
"10",
"00",
"01",
"01",
"11",
"01",
"10",
"11",
"00",
"00",
"01",
"10",
"10",
"11",
"00",
"00",
"01",
"10",
"11",
"11",
"11",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"11",
"01",
"01",
"01",
"00",
"11",
"01",
"01",
"00",
"00",
"01",
"01",
"11",
"10",
"01",
"01",
"01",
"10",
"01",
"11",
"10",
"01",
"11",
"11",
"00",
"01",
"11",
"00",
"11",
"00",
"10",
"11",
"00",
"11",
"00",
"10",
"11",
"11",
"00",
"10",
"11",
"01",
"01",
"01",
"00",
"01",
"01",
"01",
"10",
"01",
"01",
"10",
"11",
"11",
"10",
"11",
"11",
"01",
"01",
"10",
"10",
"10",
"10",
"11",
"01",
"01",
"11",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"00",
"00",
"01",
"11",
"10",
"11",
"01",
"10",
"00",
"10",
"01",
"10",
"00",
"00",
"01",
"11",
"10",
"00",
"11",
"00",
"11",
"01",
"00",
"10",
"00",
"00",
"01",
"01",
"00",
"10",
"10",
"01",
"11",
"01",
"00",
"01",
"10",
"11",
"10",
"00",
"01",
"00",
"11",
"11",
"10",
"10",
"10",
"00",
"00",
"01",
"11",
"11",
"10",
"01",
"11",
"01",
"01",
"11",
"10",
"00",
"11",
"00",
"10",
"11",
"01",
"10",
"11",
"11",
"01",
"00",
"10",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"01",
"11",
"00",
"00",
"01",
"10",
"01",
"11",
"11",
"11",
"11",
"01",
"10",
"01",
"10",
"00",
"01",
"10",
"10",
"11",
"01",
"01",
"01",
"10",
"10",
"10",
"11",
"11",
"00",
"11",
"10",
"00",
"01",
"01",
"11",
"00",
"01",
"01",
"01",
"00",
"11",
"10",
"10",
"01",
"10",
"10",
"11",
"11",
"00",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"01",
"01",
"11",
"10",
"00",
"10",
"10",
"10",
"00",
"10",
"11",
"00",
"11",
"10",
"10",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"11",
"11",
"11",
"11",
"11",
"11",
"00",
"11",
"00",
"11",
"01",
"01",
"00",
"01",
"01",
"00",
"00",
"00",
"10",
"01",
"11",
"11",
"01",
"10",
"00",
"10",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"10",
"10",
"10",
"10",
"10",
"10",
"01",
"00",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"00",
"00",
"10",
"10",
"00",
"01",
"01",
"00",
"00",
"01",
"10",
"00",
"10",
"10",
"11",
"10",
"11",
"00",
"01",
"10",
"11",
"00",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"01",
"01",
"00",
"01",
"10",
"00",
"01",
"10",
"01",
"10",
"00",
"01",
"01",
"01",
"10",
"11",
"10",
"10",
"10",
"10",
"00",
"01",
"10",
"10",
"00",
"01",
"11",
"10",
"00",
"00",
"00",
"00",
"11",
"00",
"10",
"11",
"11",
"11",
"11",
"00",
"11",
"10",
"01",
"11",
"11",
"10",
"10",
"01",
"10",
"01",
"10",
"01",
"10",
"00",
"11",
"01",
"10",
"11",
"00",
"11",
"00",
"11",
"01",
"01",
"10",
"00",
"11",
"11",
"01",
"10",
"11",
"01",
"01",
"11",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"01",
"11",
"01",
"01",
"00",
"11",
"00",
"10",
"11",
"10",
"11",
"01",
"00",
"00",
"01",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"01",
"10",
"11",
"10",
"01",
"00",
"00",
"11",
"01",
"00",
"01",
"11",
"00",
"11",
"00",
"00",
"10",
"01",
"01",
"10",
"00",
"00",
"10",
"00",
"00",
"00",
"01",
"01",
"10",
"10",
"11",
"01",
"01",
"01",
"11",
"11",
"10",
"01",
"10",
"10",
"00",
"00",
"01",
"10",
"01",
"01",
"01",
"00",
"00",
"00",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"11",
"11",
"11",
"00",
"11",
"11",
"01",
"10",
"01",
"01",
"00",
"01",
"00",
"11",
"10",
"00",
"10",
"00",
"00",
"00",
"11",
"11",
"00",
"01",
"10",
"01",
"10",
"00",
"11",
"00",
"10",
"10",
"01",
"11",
"11",
"11",
"00",
"11",
"00",
"11",
"01",
"00",
"10",
"00",
"11",
"00",
"10",
"11",
"01",
"11",
"10",
"10",
"10",
"00",
"00",
"10",
"11",
"10",
"11",
"00",
"11",
"10",
"01",
"10",
"01",
"10",
"10",
"11",
"00",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"11",
"00",
"10",
"01",
"01",
"11",
"11",
"01",
"01",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"00",
"11",
"11",
"10",
"01",
"10",
"01",
"00",
"10",
"10",
"01",
"10",
"01",
"00",
"10",
"00",
"10",
"00",
"10",
"00",
"10",
"01",
"11",
"10",
"11",
"01",
"01",
"00",
"11",
"00",
"00",
"10",
"11",
"11",
"10",
"11",
"11",
"00",
"00",
"00",
"10",
"00",
"10",
"01",
"01",
"10",
"00",
"01",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"00",
"11",
"00",
"11",
"10",
"01",
"01",
"10",
"01",
"11",
"00",
"10",
"00",
"10",
"00",
"01",
"01",
"11",
"11",
"11",
"10",
"00",
"01",
"01",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"11",
"01",
"01",
"10",
"01",
"11",
"00",
"11",
"11",
"01",
"11",
"01",
"10",
"00",
"00",
"11",
"00",
"10",
"00",
"11",
"11",
"10",
"01",
"10",
"00",
"00",
"00",
"11",
"10",
"01",
"01",
"11",
"00",
"00",
"11",
"10",
"01",
"11",
"01",
"01",
"10",
"01",
"01",
"10",
"01",
"11",
"01",
"00",
"01",
"01",
"01",
"11",
"11",
"01",
"00",
"00",
"11",
"10",
"01",
"00",
"00",
"10",
"00",
"10",
"11",
"10",
"11",
"01",
"11",
"10",
"10",
"11",
"11",
"00",
"01",
"00",
"11",
"11",
"00",
"00",
"01",
"00",
"00",
"11",
"11",
"00",
"01",
"10",
"11",
"01",
"00",
"01",
"01",
"11",
"10",
"11",
"11",
"01",
"00",
"01",
"10",
"11",
"11",
"11",
"00",
"01",
"01",
"01",
"01",
"10",
"10",
"01",
"11",
"01",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"01",
"10",
"00",
"10",
"00",
"01",
"10",
"01",
"00",
"00",
"01",
"11",
"01",
"11",
"10",
"11",
"10",
"01",
"11",
"11",
"00",
"11",
"01",
"00",
"00",
"01",
"00",
"10",
"11",
"00",
"00",
"11",
"01",
"01",
"00",
"00",
"00",
"00",
"11",
"11",
"00",
"10",
"00",
"11",
"11",
"00",
"01",
"01",
"11",
"01",
"11",
"10",
"11",
"10",
"00",
"00",
"00",
"10",
"11",
"00",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"10",
"01",
"11",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"11",
"00",
"00",
"10",
"11",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"11",
"11",
"01",
"01",
"10",
"11",
"10",
"00",
"01",
"01",
"10",
"00",
"01",
"01",
"00",
"11",
"11",
"01",
"10",
"10",
"01",
"00",
"00",
"10",
"10",
"00",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"10",
"11",
"01",
"00",
"11",
"10",
"00",
"11",
"00",
"00",
"11",
"10",
"00",
"01",
"00",
"00",
"00",
"01",
"11",
"11",
"00",
"00",
"00",
"01",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"01",
"11",
"01",
"11",
"10",
"00",
"11",
"00",
"11",
"00",
"10",
"00",
"11",
"00",
"01",
"11",
"01",
"00",
"00",
"11",
"00",
"01",
"00",
"10",
"01",
"10",
"01",
"10",
"00",
"10",
"00",
"11",
"00",
"01",
"11",
"10",
"00",
"00",
"10",
"01",
"00",
"00",
"00",
"10",
"01",
"00",
"10",
"11",
"01",
"00",
"01",
"00",
"11",
"10",
"10",
"00",
"01",
"10",
"10",
"00",
"00",
"01",
"10",
"00",
"01",
"10",
"00",
"11",
"00",
"11",
"11",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"00",
"00",
"11",
"01",
"00",
"00",
"11",
"10",
"00",
"11",
"00",
"11",
"10",
"01",
"01",
"00",
"01",
"10",
"00",
"11",
"11",
"10",
"10",
"00",
"01",
"00",
"01",
"00",
"00",
"01",
"10",
"10",
"01",
"01",
"11",
"11",
"00",
"10",
"00",
"11",
"10",
"10",
"01",
"10",
"01",
"11",
"01",
"11",
"00",
"11",
"01",
"10",
"00",
"00",
"10",
"01",
"01",
"11",
"11",
"01",
"00",
"11",
"00",
"00",
"10",
"11",
"10",
"11",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"01",
"01",
"01",
"11",
"10",
"10",
"01",
"00",
"10",
"11",
"00",
"10",
"01",
"00",
"10",
"01",
"11",
"11",
"00",
"01",
"00",
"00",
"11",
"00",
"10",
"10",
"11",
"11",
"10",
"10",
"11",
"01",
"10",
"00",
"00",
"10",
"11",
"01",
"00",
"11",
"11",
"11",
"10",
"00",
"00",
"10",
"00",
"01",
"11",
"10",
"01",
"11",
"11",
"10",
"00",
"10",
"00",
"00",
"01",
"10",
"11",
"10",
"01",
"10",
"00",
"10",
"11",
"01",
"11",
"10",
"00",
"10",
"11",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"11",
"01",
"01",
"10",
"11",
"11",
"01",
"10",
"11",
"01",
"10",
"00",
"10",
"11",
"00",
"01",
"01",
"00",
"01",
"00",
"01",
"01",
"00",
"11",
"01",
"10",
"00",
"00",
"00",
"11",
"10",
"00",
"10",
"11",
"00",
"00",
"01",
"11",
"00",
"00",
"00",
"11",
"00",
"00",
"10",
"10",
"01",
"01",
"00",
"11",
"01",
"10",
"01",
"11",
"11",
"00",
"10",
"10",
"00",
"00",
"11",
"00",
"10",
"00",
"00",
"11",
"01",
"00",
"11",
"00",
"01",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"00",
"11",
"10",
"10",
"00",
"10",
"00",
"10",
"11",
"11",
"01",
"10",
"01",
"11",
"00",
"00",
"00",
"01",
"01",
"01",
"10",
"00",
"00",
"11",
"10",
"11",
"01",
"10",
"00",
"11",
"11",
"10",
"10",
"10",
"00",
"11",
"00",
"10",
"00",
"10",
"01",
"10",
"01",
"10",
"10",
"01",
"01",
"11",
"00",
"11",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"01",
"10",
"10",
"00",
"10",
"01",
"11",
"00",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"10",
"00",
"01",
"00",
"11",
"10",
"10",
"10",
"00",
"00",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"10",
"10",
"10",
"01",
"11",
"01",
"00",
"10",
"11",
"10",
"00",
"00",
"10",
"11",
"01",
"10",
"10",
"00",
"01",
"11",
"01",
"00",
"00",
"10",
"11",
"01",
"00",
"11",
"01",
"01",
"10",
"11",
"00",
"10",
"00",
"01",
"10",
"00",
"10",
"10",
"10",
"00",
"11",
"11",
"11",
"00",
"11",
"11",
"01",
"00",
"01",
"11",
"10",
"01",
"11",
"10",
"01",
"01",
"11",
"00",
"10",
"11",
"01",
"00",
"10",
"01",
"01",
"01",
"00",
"01",
"00",
"01",
"11",
"00",
"01",
"10",
"10",
"01",
"11",
"10",
"00",
"01",
"10",
"01",
"00",
"00",
"10",
"00",
"00",
"11",
"11",
"00",
"01",
"00",
"11",
"10",
"11",
"11",
"00",
"10",
"10",
"10",
"01",
"01",
"00",
"11",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"01",
"10",
"00",
"10",
"11",
"10",
"11",
"01",
"00",
"01",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"00",
"01",
"10",
"10",
"00",
"11",
"10",
"01",
"01",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"10",
"10",
"11",
"10",
"01",
"01",
"10",
"10",
"00",
"00",
"00",
"11",
"10",
"10",
"10",
"00",
"11",
"10",
"00",
"11",
"11",
"00",
"01",
"10",
"00",
"01",
"10",
"00",
"11",
"11",
"00",
"00",
"11",
"11",
"10",
"10",
"01",
"10",
"10",
"10",
"11",
"10",
"00",
"11",
"11",
"00",
"11",
"10",
"00",
"11",
"01",
"11",
"11",
"00",
"11",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"11",
"11",
"00",
"10",
"00",
"00",
"01",
"10",
"10",
"11",
"10",
"11",
"00",
"10",
"11",
"01",
"10",
"11",
"11",
"11",
"00",
"11",
"00",
"10",
"01",
"11",
"00",
"10",
"01",
"10",
"01",
"10",
"11",
"01",
"00",
"00",
"01",
"11",
"00",
"01",
"01",
"00",
"11",
"11",
"10",
"00",
"01",
"01",
"10",
"00",
"11",
"10",
"11",
"00",
"10",
"10",
"10",
"11",
"00",
"00",
"11",
"10",
"11",
"00",
"01",
"01",
"11",
"01",
"01",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"01",
"10",
"10",
"10",
"11",
"00",
"01",
"10",
"11",
"10",
"01",
"11",
"01",
"01",
"11",
"11",
"00",
"11",
"00",
"11",
"11",
"00",
"11",
"11",
"10",
"01",
"00",
"00",
"11",
"00",
"00",
"11",
"01",
"00",
"01",
"00",
"10",
"01",
"10",
"11",
"10",
"10",
"00",
"11",
"11",
"01",
"11",
"00",
"01",
"01",
"11",
"11",
"00",
"01",
"01",
"11",
"10",
"00",
"10",
"11",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"11",
"00",
"01",
"11",
"10",
"11",
"00",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"01",
"00",
"10",
"10",
"00",
"01",
"10",
"00",
"10",
"00",
"00",
"01",
"00",
"00",
"00",
"01",
"01",
"11",
"11",
"10",
"11",
"01",
"11",
"11",
"11",
"11",
"01",
"10",
"11",
"00",
"00",
"11",
"10",
"00",
"11",
"11",
"11",
"11",
"00",
"00",
"10",
"01",
"01",
"11",
"00",
"10",
"11",
"11",
"00",
"00",
"00",
"11",
"11",
"00",
"10",
"01",
"01",
"11",
"00",
"01",
"01",
"11",
"00",
"00",
"10",
"00",
"11",
"00",
"01",
"00",
"10",
"01",
"00",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"00",
"11",
"00",
"10",
"11",
"10",
"01",
"00",
"01",
"11",
"01",
"10",
"00",
"00",
"11",
"00",
"11",
"01",
"10",
"10",
"10",
"10",
"01",
"01",
"11",
"11",
"11",
"10",
"11",
"11",
"11",
"10",
"00",
"00",
"01",
"10",
"10",
"11",
"10",
"11",
"10",
"11",
"10",
"00",
"01",
"01",
"01",
"11",
"11",
"00",
"00",
"00",
"11",
"00",
"11",
"10",
"00",
"11",
"01",
"10",
"00",
"00",
"00",
"01",
"10",
"00",
"11",
"00",
"11",
"11",
"00",
"10",
"11",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"01",
"01",
"10",
"01",
"11",
"01",
"01",
"11",
"11",
"11",
"01",
"11",
"10",
"00",
"10",
"11",
"00",
"01",
"11",
"01",
"10",
"00",
"11",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"10",
"01",
"10",
"11",
"00",
"11",
"10",
"11",
"00",
"01",
"11",
"10",
"00",
"11",
"01",
"01",
"00",
"10",
"01",
"00",
"10",
"00",
"00",
"01",
"01",
"00",
"01",
"01",
"01",
"01",
"00",
"10",
"11",
"00",
"00",
"01",
"11",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"00",
"00",
"11",
"11",
"01",
"10",
"11",
"01",
"00",
"10",
"01",
"10",
"10",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"10",
"11",
"11",
"00",
"00",
"11",
"11",
"00",
"00",
"11",
"10",
"11",
"11",
"00",
"00",
"11",
"00",
"01",
"10",
"00",
"10",
"00",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"01",
"10",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"01",
"00",
"11",
"10",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"01",
"11",
"01",
"01",
"10",
"10",
"00",
"11",
"11",
"10",
"00",
"01",
"11",
"01",
"00",
"11",
"11",
"01",
"00",
"01",
"11",
"10",
"10",
"00",
"01",
"01",
"10",
"10",
"11",
"11",
"01",
"11",
"00",
"00",
"00",
"01",
"10",
"11",
"10",
"00",
"00",
"11",
"00",
"10",
"00",
"10",
"01",
"11",
"01",
"10",
"00",
"11",
"00",
"01",
"11",
"11",
"01",
"01",
"11",
"01",
"11",
"01",
"01",
"10",
"10",
"00",
"11",
"10",
"01",
"11",
"10",
"10",
"00",
"11",
"11",
"10",
"11",
"01",
"00",
"10",
"01",
"00",
"00",
"01",
"10",
"01",
"00",
"01",
"10",
"00",
"01",
"11",
"11",
"11",
"11",
"01",
"01",
"11",
"00",
"11",
"11",
"01",
"10",
"11",
"01",
"10",
"00",
"11",
"10",
"11",
"10",
"01",
"00",
"10",
"10",
"10",
"11",
"00",
"01",
"11",
"11",
"11",
"00",
"00",
"00",
"01",
"01",
"00",
"10",
"01",
"11",
"10",
"00",
"01",
"10",
"10",
"00",
"01",
"11",
"00",
"01",
"10",
"00",
"00",
"10",
"10",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"11",
"00",
"10",
"01",
"11",
"01",
"10",
"01",
"10",
"11",
"01",
"01",
"00",
"01",
"00",
"01",
"11",
"10",
"00",
"00",
"10",
"01",
"11",
"00",
"11",
"01",
"01",
"10",
"00",
"11",
"11",
"11",
"10",
"01",
"11",
"00",
"10",
"11",
"00",
"10",
"01",
"01",
"00",
"01",
"11",
"11",
"00",
"10",
"00",
"10",
"00",
"10",
"00",
"01",
"10",
"01",
"11",
"11",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"11",
"10",
"01",
"01",
"01",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"00",
"10",
"00",
"10",
"00",
"10",
"10",
"10",
"01",
"01",
"11",
"10",
"11",
"10",
"10",
"10",
"11",
"01",
"11",
"10",
"10",
"00",
"01",
"10",
"11",
"01",
"00",
"11",
"10",
"10",
"00",
"11",
"10",
"01",
"01",
"00",
"00",
"01",
"01",
"01",
"01",
"11",
"00",
"10",
"01",
"10",
"10",
"11",
"11",
"01",
"10",
"00",
"10",
"10",
"00",
"01",
"10",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"11",
"10",
"01",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"10",
"11",
"00",
"10",
"11",
"01",
"00",
"10",
"10",
"11",
"11",
"00",
"11",
"00",
"11",
"01",
"00",
"11",
"11",
"00",
"10",
"01",
"00",
"10",
"10",
"01",
"11",
"01",
"10",
"10",
"10",
"11",
"11",
"11",
"10",
"11",
"10",
"10",
"10",
"00",
"10",
"10",
"01",
"10",
"10",
"00",
"01",
"10",
"10",
"00",
"11",
"11",
"01",
"11",
"01",
"00",
"10",
"00",
"00",
"11",
"01",
"00",
"00",
"10",
"11",
"01",
"01",
"01",
"01",
"10",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"10",
"00",
"00",
"10",
"00",
"01",
"11",
"01",
"11",
"00",
"10",
"11",
"01",
"11",
"11",
"01",
"00",
"01",
"11",
"01",
"10",
"10",
"11",
"10",
"00",
"11",
"00",
"10",
"10",
"01",
"10",
"00",
"10",
"00",
"00",
"11",
"01",
"00",
"10",
"00",
"11",
"01",
"00",
"10",
"01",
"11",
"11",
"00",
"11",
"01",
"10",
"10",
"01",
"01",
"00",
"01",
"01",
"01",
"10",
"01",
"00",
"10",
"00",
"10",
"11",
"11",
"11",
"10",
"00",
"10",
"11",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"00",
"00",
"10",
"00",
"10",
"10",
"01",
"00",
"01",
"11",
"00",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"10",
"01",
"01",
"00",
"11",
"11",
"01",
"01",
"01",
"01",
"00",
"11",
"01",
"10",
"01",
"11",
"10",
"01",
"10",
"01",
"00",
"11",
"11",
"11",
"01",
"00",
"10",
"01",
"11",
"11",
"10",
"10",
"10",
"00",
"00",
"11",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"00",
"00",
"00",
"10",
"10",
"01",
"10",
"00",
"00",
"10",
"10",
"11",
"01",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"11",
"10",
"10",
"10",
"10",
"10",
"01",
"11",
"00",
"01",
"01",
"01",
"10",
"01",
"00",
"00",
"01",
"00",
"00",
"11",
"11",
"10",
"11",
"11",
"10",
"01",
"10",
"11",
"00",
"00",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"11",
"10",
"10",
"11",
"11",
"00",
"01",
"11",
"00",
"01",
"11",
"00",
"01",
"01",
"00",
"11",
"10",
"00",
"00",
"01",
"00",
"00",
"01",
"01",
"00",
"10",
"01",
"11",
"01",
"01",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"10",
"10",
"11",
"11",
"00",
"10",
"11",
"11",
"00",
"10",
"01",
"11",
"10",
"01",
"01",
"00",
"10",
"00",
"11",
"11",
"11",
"11",
"00",
"00",
"01",
"00",
"10",
"11",
"01",
"10",
"11",
"10",
"10",
"01",
"11",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"01",
"11",
"11",
"10",
"11",
"11",
"01",
"00",
"00",
"00",
"00",
"11",
"11",
"10",
"11",
"01",
"00",
"01",
"10",
"01",
"01",
"10",
"10",
"00",
"11",
"01",
"11",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"00",
"00",
"01",
"00",
"11",
"11",
"10",
"01",
"01",
"10",
"10",
"01",
"00",
"00",
"00",
"00",
"11",
"00",
"01",
"10",
"10",
"01",
"01",
"00",
"11",
"11",
"10",
"11",
"10",
"00",
"00",
"00",
"01",
"11",
"11",
"01",
"01",
"00",
"11",
"00",
"00",
"10",
"01",
"11",
"01",
"01",
"10",
"00",
"01",
"00",
"00",
"00",
"01",
"01",
"00",
"10",
"11",
"11",
"11",
"01",
"11",
"01",
"00",
"01",
"00",
"11",
"11",
"10",
"11",
"01",
"01",
"10",
"10",
"01",
"00",
"00",
"10",
"10",
"10",
"01",
"00",
"00",
"11",
"01",
"00",
"00",
"00",
"01",
"11",
"01",
"11",
"01",
"10",
"11",
"00",
"01",
"11",
"11",
"10",
"00",
"10",
"00",
"00",
"10",
"00",
"00",
"10",
"01",
"00",
"10",
"00",
"10",
"01",
"10",
"01",
"00",
"00",
"11",
"00",
"11",
"01",
"11",
"00",
"01",
"11",
"01",
"11",
"00",
"01",
"10",
"01",
"01",
"01",
"00",
"11",
"00",
"00",
"01",
"01",
"11",
"11",
"11",
"10",
"00",
"10",
"01",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"01",
"00",
"00",
"10",
"11",
"10",
"10",
"10",
"00",
"10",
"11",
"00",
"01",
"00",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"01",
"11",
"10",
"11",
"00",
"00",
"10",
"00",
"11",
"10",
"01",
"10",
"11",
"01",
"11",
"10",
"00",
"11",
"10",
"10",
"00",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"00",
"00",
"00",
"01",
"10",
"10",
"11",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"11",
"11",
"11",
"00",
"10",
"11",
"10",
"10",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"01",
"01",
"11",
"00",
"01",
"00",
"10",
"10",
"10",
"11",
"00",
"11",
"11",
"01",
"11",
"01",
"01",
"00",
"01",
"10",
"11",
"01",
"11",
"00",
"01",
"01",
"11",
"10",
"10",
"11",
"10",
"00",
"00",
"01",
"10",
"10",
"01",
"00",
"01",
"00",
"00",
"00",
"11",
"10",
"00",
"10",
"00",
"01",
"01",
"11",
"01",
"11",
"00",
"01",
"11",
"10",
"10",
"10",
"01",
"00",
"10",
"10",
"01",
"01",
"10",
"00",
"11",
"00",
"00",
"11",
"00",
"00",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"01",
"00",
"11",
"01",
"01",
"00",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"00",
"00",
"10",
"11",
"10",
"00",
"11",
"11",
"10",
"01",
"10",
"11",
"01",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"01",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"00",
"11",
"10",
"00",
"10",
"11",
"01",
"11",
"11",
"01",
"00",
"11",
"10",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"01",
"11",
"10",
"00",
"00",
"01",
"10",
"11",
"01",
"10",
"10",
"10",
"10",
"01",
"01",
"11",
"01",
"01",
"00",
"00",
"00",
"00",
"01",
"01",
"10",
"11",
"10",
"01",
"00",
"00",
"01",
"01",
"01",
"01",
"11",
"00",
"10",
"10",
"00",
"10",
"11",
"11",
"11",
"10",
"10",
"11",
"10",
"10",
"00",
"11",
"10",
"11",
"00",
"01",
"01",
"01",
"00",
"11",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"11",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"01",
"11",
"01",
"01",
"00",
"10",
"00",
"01",
"00",
"01",
"00",
"00",
"11",
"11",
"10",
"01",
"11",
"11",
"01",
"10",
"01",
"00",
"00",
"01",
"11",
"00",
"01",
"01",
"10",
"01",
"01",
"11",
"11",
"01",
"11",
"01",
"01",
"10",
"01",
"10",
"10",
"00",
"00",
"11",
"10",
"01",
"01",
"11",
"00",
"01",
"10",
"11",
"11",
"11",
"10",
"11",
"11",
"01",
"10",
"11",
"00",
"10",
"01",
"01",
"00",
"01",
"00",
"10",
"10",
"10",
"10",
"11",
"10",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"00",
"11",
"11",
"10",
"11",
"00",
"01",
"10",
"11",
"00",
"11",
"01",
"01",
"00",
"01",
"00",
"10",
"11",
"11",
"10",
"11",
"00",
"01",
"00",
"10",
"11",
"11",
"00",
"01",
"00",
"00",
"00",
"10",
"01",
"01",
"00",
"00",
"10",
"11",
"10",
"10",
"11",
"10",
"11",
"10",
"10",
"00",
"00",
"01",
"00",
"01",
"11",
"01",
"01",
"10",
"10",
"11",
"00",
"00",
"11",
"11",
"10",
"10",
"11",
"01",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"00",
"01",
"11",
"10",
"01",
"10",
"10",
"11",
"10",
"10",
"01",
"10",
"01",
"00",
"01",
"00",
"11",
"01",
"01",
"10",
"01",
"00",
"01",
"11",
"00",
"10",
"00",
"01",
"01",
"01",
"10",
"10",
"00",
"10",
"00",
"11",
"00",
"01",
"00",
"00",
"00",
"10",
"00",
"11",
"11",
"11",
"01",
"00",
"10",
"00",
"00",
"00",
"01",
"11",
"10",
"11",
"10",
"01",
"00",
"10",
"01",
"00",
"10",
"00",
"01",
"11",
"00",
"00",
"01",
"00",
"10",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"00",
"10",
"00",
"11",
"01",
"11",
"11",
"00",
"10",
"10",
"11",
"10",
"11",
"10",
"00",
"11",
"11",
"00",
"00",
"11",
"00",
"10",
"00",
"11",
"10",
"11",
"00",
"00",
"01",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"00",
"01",
"01",
"01",
"11",
"10",
"01",
"10",
"00",
"10",
"10",
"00",
"01",
"11",
"00",
"01",
"10",
"10",
"01",
"11",
"00",
"01",
"00",
"00",
"11",
"11",
"10",
"11",
"00",
"11",
"01",
"01",
"00",
"10",
"01",
"11",
"10",
"01",
"00",
"11",
"10",
"11",
"01",
"00",
"11",
"10",
"10",
"11",
"00",
"01",
"00",
"10",
"11",
"10",
"01",
"00",
"10",
"10",
"10",
"10",
"11",
"00",
"00",
"10",
"11",
"01",
"10",
"10",
"00",
"00",
"00",
"10",
"10",
"00",
"10",
"11",
"00",
"10",
"00",
"10",
"10",
"01",
"11",
"11",
"00",
"00",
"00",
"01",
"10",
"00",
"10",
"11",
"11",
"10",
"01",
"01",
"01",
"10",
"01",
"11",
"11",
"10",
"00",
"00",
"00",
"10",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"00",
"00",
"00",
"01",
"11",
"11",
"00",
"11",
"00",
"01",
"01",
"11",
"00",
"11",
"01",
"10",
"10",
"11",
"10",
"11",
"01",
"10",
"11",
"00",
"01",
"10",
"11",
"00",
"10",
"00",
"11",
"00",
"11",
"00",
"01",
"11",
"10",
"01",
"01",
"11",
"11",
"11",
"01",
"11",
"11",
"00",
"00",
"00",
"11",
"10",
"11",
"00",
"00",
"00",
"10",
"11",
"01",
"11",
"01",
"00",
"01",
"01",
"10",
"11",
"01",
"11",
"00",
"11",
"01",
"10",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"11",
"00",
"00",
"01",
"00",
"00",
"10",
"01",
"11",
"10",
"00",
"11",
"01",
"00",
"11",
"11",
"10",
"10",
"11",
"01",
"10",
"11",
"11",
"00",
"10",
"10",
"10",
"10",
"00",
"01",
"10",
"11",
"01",
"10",
"10",
"01",
"00",
"00",
"11",
"11",
"01",
"11",
"10",
"01",
"10",
"01",
"11",
"10",
"11",
"11",
"11",
"01",
"11",
"10",
"01",
"01",
"00",
"01",
"10",
"11",
"01",
"01",
"00",
"10",
"01",
"11",
"01",
"00",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"11",
"00",
"11",
"00",
"11",
"10",
"00",
"00",
"11",
"00",
"00",
"01",
"11",
"00",
"10",
"00",
"10",
"11",
"01",
"01",
"11",
"10",
"11",
"10",
"01",
"11",
"01",
"11",
"00",
"11",
"00",
"01",
"11",
"10",
"01",
"11",
"01",
"00",
"01",
"10",
"00",
"00",
"11",
"01",
"11",
"00",
"11",
"01",
"10",
"00",
"00",
"01",
"11",
"11",
"01",
"10",
"11",
"10",
"01",
"00",
"01",
"00",
"00",
"10",
"11",
"10",
"01",
"10",
"11",
"10",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"10",
"11",
"00",
"10",
"01",
"00",
"10",
"10",
"01",
"01",
"01",
"11",
"11",
"10",
"11",
"11",
"01",
"01",
"01",
"00",
"00",
"10",
"10",
"00",
"00",
"11",
"00",
"11",
"00",
"10",
"00",
"01",
"01",
"11",
"00",
"10",
"11",
"00",
"11",
"10",
"11",
"00",
"11",
"10",
"11",
"10",
"01",
"00",
"01",
"11",
"01",
"11",
"10",
"00",
"10",
"01",
"11",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"10",
"10",
"10",
"10",
"11",
"11",
"10",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"00",
"01",
"11",
"00",
"00",
"11",
"01",
"00",
"00",
"00",
"11",
"10",
"00",
"01",
"01",
"10",
"01",
"00",
"11",
"11",
"10",
"00",
"01",
"11",
"01",
"10",
"00",
"01",
"00",
"11",
"00",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"00",
"01",
"10",
"10",
"00",
"00",
"10",
"01",
"10",
"00",
"11",
"11",
"11",
"00",
"11",
"10",
"00",
"00",
"11",
"00",
"10",
"10",
"00",
"00",
"10",
"10",
"00",
"00",
"11",
"00",
"11",
"00",
"10",
"01",
"11",
"11",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"00",
"10",
"01",
"11",
"01",
"01",
"00",
"11",
"10",
"11",
"00",
"11",
"01",
"11",
"00",
"11",
"10",
"11",
"10",
"11",
"00",
"10",
"01",
"11",
"10",
"11",
"01",
"00",
"00",
"01",
"11",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"00",
"11",
"11",
"00",
"01",
"01",
"00",
"11",
"10",
"00",
"00",
"10",
"01",
"11",
"00",
"01",
"11",
"01",
"00",
"11",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"00",
"00",
"10",
"01",
"10",
"01",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"10",
"01",
"00",
"11",
"10",
"00",
"01",
"01",
"00",
"11",
"10",
"00",
"10",
"11",
"00",
"01",
"11",
"00",
"11",
"00",
"11",
"10",
"00",
"00",
"01",
"01",
"11",
"00",
"00",
"10",
"10",
"00",
"11",
"01",
"11",
"00",
"00",
"01",
"01",
"10",
"11",
"10",
"01",
"01",
"11",
"01",
"10",
"11",
"11",
"11",
"01",
"11",
"00",
"11",
"10",
"11",
"11",
"10",
"00",
"01",
"01",
"00",
"11",
"00",
"11",
"10",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"01",
"10",
"11",
"00",
"10",
"01",
"10",
"10",
"00",
"11",
"01",
"10",
"01",
"10",
"00",
"01",
"01",
"11",
"11",
"00",
"00",
"01",
"11",
"10",
"00",
"00",
"11",
"11",
"01",
"01",
"10",
"01",
"11",
"10",
"10",
"11",
"01",
"10",
"10",
"11",
"01",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"11",
"10",
"01",
"00",
"00",
"10",
"01",
"10",
"10",
"00",
"10",
"00",
"11",
"11",
"01",
"01",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"11",
"10",
"10",
"10",
"00",
"01",
"10",
"00",
"01",
"11",
"11",
"11",
"00",
"11",
"11",
"10",
"01",
"10",
"10",
"11",
"11",
"10",
"01",
"01",
"01",
"11",
"11",
"11",
"01",
"10",
"00",
"10",
"00",
"11",
"00",
"01",
"01",
"11",
"10",
"10",
"00",
"10",
"10",
"01",
"10",
"01",
"11",
"11",
"11",
"11",
"01",
"10",
"01",
"10",
"01",
"01",
"00",
"10",
"01",
"11",
"01",
"01",
"00",
"01",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"00",
"10",
"00",
"10",
"10",
"10",
"10",
"10",
"10",
"00",
"11",
"10",
"01",
"00",
"00",
"01",
"10",
"01",
"10",
"11",
"10",
"01",
"01",
"10",
"11",
"00",
"00",
"11",
"00",
"01",
"01",
"00",
"00",
"01",
"11",
"11",
"11",
"00",
"11",
"10",
"10",
"01",
"11",
"11",
"11",
"10",
"00",
"10",
"11",
"00",
"11",
"00",
"11",
"10",
"10",
"11",
"00",
"01",
"11",
"11",
"01",
"00",
"01",
"01",
"00",
"11",
"10",
"11",
"10",
"01",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"01",
"10",
"01",
"00",
"10",
"00",
"10",
"01",
"01",
"11",
"01",
"11",
"10",
"01",
"01",
"01",
"01",
"10",
"01",
"11",
"11",
"00",
"11",
"11",
"11",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"00",
"01",
"01",
"10",
"10",
"11",
"00",
"01",
"01",
"10",
"10",
"10",
"01",
"00",
"00",
"01",
"00",
"00",
"11",
"11",
"11",
"01",
"11",
"00",
"00",
"10",
"01",
"01",
"10",
"00",
"00",
"00",
"10",
"01",
"11",
"10",
"10",
"10",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"00",
"11",
"00",
"11",
"10",
"01",
"01",
"00",
"00",
"01",
"11",
"00",
"00",
"01",
"01",
"00",
"01",
"10",
"10",
"10",
"10",
"11",
"00",
"11",
"11",
"10",
"11",
"10",
"00",
"01",
"10",
"01",
"10",
"11",
"01",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"01",
"00",
"01",
"00",
"00",
"00",
"01",
"00",
"01",
"00",
"00",
"10",
"10",
"11",
"11",
"00",
"00",
"10",
"00",
"00",
"11",
"00",
"10",
"00",
"11",
"01",
"11",
"01",
"10",
"00",
"01",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"01",
"01",
"01",
"00",
"01",
"10",
"10",
"10",
"11",
"11",
"00",
"01",
"00",
"01",
"11",
"01",
"01",
"11",
"10",
"11",
"10",
"11",
"11",
"11",
"11",
"00",
"01",
"00",
"11",
"00",
"10",
"10",
"11",
"00",
"00",
"10",
"10",
"01",
"11",
"01",
"01",
"11",
"00",
"01",
"00",
"10",
"00",
"10",
"11",
"00",
"11",
"11",
"00",
"00",
"10",
"01",
"10",
"11",
"01",
"10",
"10",
"01",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"10",
"00",
"01",
"11",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"10",
"00",
"11",
"10",
"01",
"00",
"11",
"00",
"01",
"11",
"01",
"01",
"00",
"11",
"11",
"10",
"01",
"10",
"00",
"11",
"10",
"00",
"00",
"10",
"00",
"10",
"10",
"00",
"11",
"00",
"10",
"11",
"11",
"11",
"01",
"10",
"01",
"00",
"00",
"00",
"11",
"10",
"00",
"11",
"10",
"01",
"11",
"11",
"00",
"11",
"10",
"11",
"11",
"11",
"11",
"11",
"10",
"00",
"00",
"01",
"00",
"10",
"01",
"01",
"01",
"01",
"10",
"01",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"11",
"00",
"11",
"00",
"00",
"10",
"11",
"01",
"00",
"10",
"10",
"01",
"00",
"10",
"11",
"10",
"00",
"01",
"11",
"00",
"01",
"01",
"11",
"10",
"11",
"10",
"01",
"10",
"00",
"10",
"11",
"10",
"01",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"10",
"00",
"01",
"11",
"00",
"01",
"00",
"00",
"10",
"11",
"10",
"00",
"10",
"00",
"10",
"00",
"01",
"01",
"11",
"00",
"10",
"10",
"10",
"10",
"00",
"00",
"10",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"00",
"11",
"00",
"10",
"01",
"00",
"01",
"00",
"00",
"11",
"11",
"00",
"10",
"10",
"00",
"01",
"10",
"11",
"00",
"10",
"11",
"00",
"10",
"11",
"11",
"00",
"11",
"01",
"00",
"00",
"11",
"00",
"10",
"01",
"00",
"00",
"11",
"01",
"11",
"00",
"01",
"00",
"01",
"10",
"11",
"00",
"11",
"00",
"11",
"11",
"10",
"10",
"00",
"00",
"01",
"01",
"01",
"10",
"11",
"11",
"10",
"10",
"00",
"01",
"10",
"00",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"01",
"10",
"10",
"10",
"11",
"01",
"10",
"10",
"10",
"01",
"11",
"01",
"10",
"00",
"00",
"11",
"01",
"01",
"11",
"10",
"00",
"11",
"10",
"00",
"11",
"01",
"01",
"11",
"01",
"01",
"10",
"11",
"10",
"00",
"11",
"10",
"00",
"10",
"10",
"00",
"00",
"00",
"00",
"11",
"01",
"10",
"01",
"00",
"00",
"00",
"00",
"10",
"01",
"10",
"00",
"01",
"00",
"01",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"01",
"11",
"11",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"10",
"00",
"11",
"11",
"00",
"11",
"01",
"00",
"01",
"00",
"11",
"01",
"01",
"10",
"11",
"01",
"01",
"11",
"00",
"10",
"00",
"10",
"01",
"11",
"10",
"01",
"11",
"11",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"00",
"10",
"00",
"11",
"01",
"10",
"11",
"11",
"00",
"01",
"01",
"10",
"00",
"01",
"01",
"00",
"10",
"01",
"11",
"01",
"11",
"00",
"00",
"10",
"10",
"10",
"11",
"11",
"01",
"10",
"10",
"10",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"10",
"11",
"11",
"00",
"11",
"00",
"00",
"10",
"10",
"00",
"01",
"00",
"01",
"10",
"10",
"10",
"01",
"00",
"01",
"01",
"10",
"01",
"00",
"00",
"10",
"00",
"10",
"10",
"11",
"01",
"00",
"01",
"00",
"10",
"10",
"00",
"10",
"00",
"01",
"01",
"01",
"00",
"10",
"01",
"00",
"11",
"10",
"10",
"01",
"01",
"00",
"10",
"11",
"01",
"11",
"00",
"11",
"01",
"00",
"01",
"01",
"11",
"01",
"11",
"10",
"11",
"11",
"10",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"10",
"10",
"01",
"11",
"10",
"01",
"00",
"11",
"10",
"01",
"11",
"10",
"01",
"11",
"00",
"11",
"01",
"00",
"11",
"01",
"10",
"10",
"01",
"10",
"00",
"10",
"11",
"10",
"00",
"01",
"10",
"01",
"01",
"01",
"01",
"00",
"00",
"00",
"00",
"11",
"11",
"11",
"00",
"01",
"01",
"01",
"10",
"11",
"00",
"00",
"00",
"10",
"11",
"00",
"01",
"00",
"11",
"01",
"00",
"11",
"00",
"10",
"00",
"10",
"11",
"11",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"10",
"10",
"10",
"10",
"11",
"10",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"00",
"01",
"10",
"10",
"10",
"11",
"10",
"10",
"11",
"00",
"01",
"00",
"11",
"11",
"11",
"10",
"10",
"11",
"01",
"01",
"00",
"10",
"01",
"01",
"10",
"00",
"00",
"11",
"00",
"00",
"01",
"00",
"11",
"01",
"10",
"11",
"00",
"10",
"00",
"11",
"01",
"01",
"11",
"01",
"11",
"01",
"00",
"11",
"00",
"00",
"01",
"10",
"01",
"10",
"00",
"10",
"10",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"11",
"10",
"10",
"01",
"01",
"01",
"11",
"10",
"01",
"00",
"10",
"00",
"01",
"11",
"11",
"10",
"11",
"01",
"00",
"10",
"00",
"11",
"11",
"01",
"01",
"01",
"10",
"00",
"01",
"11",
"01",
"11",
"01",
"11",
"00",
"10",
"01",
"10",
"01",
"00",
"01",
"10",
"01",
"10",
"10",
"00",
"10",
"01",
"10",
"00",
"00",
"10",
"11",
"00",
"11",
"01",
"10",
"10",
"10",
"10",
"11",
"10",
"00",
"00",
"00",
"01",
"11",
"10",
"00",
"11",
"10",
"00",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"00",
"11",
"11",
"10",
"10",
"01",
"11",
"00",
"10",
"01",
"01",
"00",
"00",
"00",
"11",
"01",
"01",
"10",
"01",
"10",
"10",
"01",
"01",
"11",
"00",
"11",
"00",
"10",
"11",
"01",
"00",
"11",
"10",
"11",
"11",
"01",
"00",
"00",
"00",
"11",
"11",
"11",
"10",
"00",
"11",
"10",
"11",
"10",
"01",
"01",
"00",
"00",
"01",
"01",
"01",
"01",
"10",
"10",
"00",
"00",
"00",
"10",
"11",
"00",
"01",
"00",
"00",
"01",
"10",
"11",
"10",
"11",
"00",
"01",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"01",
"01",
"01",
"01",
"11",
"10",
"10",
"11",
"10",
"10",
"01",
"11",
"11",
"00",
"00",
"11",
"11",
"00",
"00",
"11",
"00",
"01",
"11",
"11",
"10",
"01",
"11",
"00",
"00",
"10",
"00",
"11",
"10",
"00",
"01",
"00",
"11",
"00",
"11",
"10",
"01",
"11",
"11",
"00",
"11",
"00",
"11",
"01",
"01",
"10",
"00",
"11",
"10",
"10",
"01",
"10",
"00",
"00",
"10",
"10",
"01",
"00",
"01",
"11",
"00",
"10",
"10",
"00",
"11",
"11",
"10",
"01",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"00",
"00",
"01",
"11",
"01",
"00",
"10",
"11",
"01",
"10",
"00",
"10",
"01",
"00",
"01",
"11",
"10",
"11",
"10",
"01",
"11",
"10",
"01",
"11",
"11",
"01",
"00",
"01",
"01",
"10",
"11",
"01",
"01",
"00",
"01",
"11",
"00",
"10",
"10",
"10",
"01",
"10",
"11",
"11",
"10",
"00",
"10",
"10",
"00",
"10",
"01",
"00",
"11",
"00",
"00",
"11",
"11",
"00",
"11",
"00",
"01",
"11",
"11",
"10",
"01",
"11",
"00",
"11",
"11",
"00",
"11",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"01",
"10",
"11",
"01",
"11",
"11",
"00",
"10",
"00",
"11",
"10",
"11",
"01",
"10",
"00",
"01",
"11",
"00",
"11",
"11",
"01",
"01",
"11",
"10",
"00",
"10",
"10",
"11",
"00",
"01",
"11",
"10",
"11",
"10",
"11",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"11",
"00",
"01",
"11",
"01",
"10",
"11",
"10",
"00",
"01",
"01",
"10",
"01",
"01",
"10",
"01",
"01",
"00",
"11",
"11",
"11",
"01",
"10",
"11",
"00",
"01",
"11",
"10",
"01",
"00",
"00",
"11",
"00",
"01",
"00",
"00",
"01",
"10",
"10",
"00",
"11",
"01",
"01",
"01",
"00",
"00",
"11",
"10",
"11",
"01",
"00",
"10",
"00",
"11",
"01",
"00",
"00",
"10",
"00",
"01",
"10",
"10",
"11",
"11",
"01",
"01",
"01",
"00",
"00",
"10",
"00",
"01",
"11",
"10",
"11",
"00",
"00",
"01",
"00",
"11",
"00",
"00",
"11",
"00",
"01",
"01",
"00",
"01",
"10",
"00",
"01",
"01",
"00",
"01",
"10",
"01",
"01",
"01",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"00",
"10",
"11",
"00",
"00",
"01",
"01",
"00",
"10",
"10",
"00",
"00",
"11",
"01",
"01",
"01",
"11",
"10",
"01",
"11",
"00",
"00",
"10",
"00",
"00",
"00",
"10",
"01",
"01",
"10",
"01",
"11",
"01",
"11",
"11",
"00",
"11",
"00",
"10",
"10",
"01",
"10",
"11",
"01",
"10",
"11",
"01",
"11",
"11",
"01",
"01",
"00",
"10",
"10",
"00",
"00",
"00",
"10",
"00",
"00",
"00",
"00",
"01",
"10",
"01",
"10",
"11",
"11",
"01",
"00",
"00",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"01",
"11",
"10",
"00",
"00",
"11",
"11",
"00",
"10",
"00",
"10",
"11",
"10",
"01",
"11",
"01",
"01",
"11",
"00",
"00",
"10",
"11",
"11",
"11",
"00",
"10",
"10",
"10",
"10",
"00",
"11",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"00",
"00",
"01",
"00",
"10",
"01",
"11",
"00",
"00",
"10",
"10",
"01",
"11",
"00",
"01",
"11",
"00",
"00",
"10",
"10",
"00",
"10",
"00",
"10",
"10",
"01",
"11",
"01",
"11",
"11",
"00",
"00",
"01",
"11",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"11",
"01",
"01",
"11",
"11",
"10",
"01",
"00",
"00",
"01",
"01",
"11",
"00",
"00",
"01",
"00",
"10",
"00",
"00",
"11",
"01",
"10",
"10",
"00",
"10",
"01",
"00",
"01",
"00",
"11",
"11",
"10",
"11",
"00",
"01",
"00",
"10",
"01",
"00",
"00",
"11",
"01",
"00",
"11",
"01",
"11",
"10",
"10",
"00",
"00",
"00",
"00",
"11",
"10",
"10",
"11",
"00",
"00",
"01",
"10",
"00",
"10",
"10",
"11",
"01",
"01",
"10",
"11",
"11",
"11",
"11",
"10",
"01",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"00",
"10",
"00",
"01",
"10",
"11",
"11",
"11",
"11",
"10",
"01",
"11",
"00",
"11",
"10",
"01",
"01",
"10",
"11",
"01",
"10",
"11",
"01",
"00",
"01",
"01",
"01",
"10",
"10",
"00",
"01",
"11",
"01",
"00",
"01",
"01",
"01",
"00",
"01",
"10",
"10",
"10",
"10",
"01",
"01",
"11",
"10",
"00",
"00",
"11",
"01",
"01",
"10",
"01",
"01",
"10",
"10",
"01",
"11",
"11",
"01",
"01",
"01",
"11",
"11",
"00",
"10",
"11",
"00",
"11",
"10",
"01",
"10",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"01",
"00",
"01",
"10",
"11",
"00",
"00",
"00",
"11",
"11",
"11",
"11",
"00",
"10",
"11",
"11",
"00",
"00",
"01",
"01",
"10",
"01",
"00",
"00",
"01",
"00",
"10",
"00",
"10",
"00",
"00",
"11",
"00",
"10",
"11",
"00",
"01",
"00",
"11",
"10",
"11",
"00",
"00",
"11",
"10",
"10",
"11",
"00",
"11",
"01",
"10",
"10",
"00",
"00",
"11",
"01",
"10",
"01",
"00",
"10",
"00",
"00",
"10",
"10",
"01",
"01",
"10",
"00",
"00",
"11",
"10",
"01",
"01",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"10",
"11",
"01",
"00",
"00",
"00",
"11",
"01",
"01",
"01",
"11",
"00",
"00",
"01",
"10",
"11",
"01",
"00",
"10",
"10",
"00",
"10",
"01",
"11",
"11",
"01",
"10",
"00",
"10",
"10",
"11",
"01",
"00",
"10",
"10",
"11",
"11",
"11",
"01",
"00",
"11",
"01",
"01",
"01",
"00",
"00",
"00",
"10",
"01",
"11",
"10",
"10",
"00",
"10",
"00",
"00",
"00",
"11",
"01",
"11",
"00",
"11",
"11",
"00",
"00",
"00",
"01",
"00",
"10",
"01",
"00",
"00",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"00",
"00",
"01",
"01",
"00",
"10",
"10",
"10",
"01",
"01",
"10",
"10",
"10",
"01",
"01",
"11",
"10",
"10",
"10",
"01",
"00",
"10",
"01",
"11",
"10",
"00",
"11",
"01",
"10",
"10",
"00",
"10",
"11",
"01",
"10",
"11",
"00",
"10",
"10",
"01",
"10",
"11",
"01",
"00",
"10",
"00",
"01",
"11",
"11",
"01",
"10",
"10",
"00",
"00",
"00",
"00",
"01",
"01",
"01",
"01",
"10",
"01",
"01",
"10",
"01",
"00",
"01",
"11",
"01",
"00",
"01",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"11",
"10",
"10",
"01",
"11",
"01",
"11",
"01",
"11",
"11",
"00",
"01",
"10",
"00",
"10",
"01",
"10",
"11",
"00",
"01",
"00",
"01",
"10",
"01",
"10",
"00",
"01",
"00",
"11",
"01",
"10",
"01",
"10",
"10",
"00",
"00",
"00",
"00",
"11",
"10",
"10",
"01",
"01",
"01",
"10",
"01",
"01",
"01",
"10",
"00",
"11",
"11",
"11",
"00",
"11",
"01",
"01",
"01",
"10",
"01",
"10",
"01",
"00",
"10",
"11",
"01",
"10",
"11",
"01",
"11",
"00",
"00",
"00",
"10",
"11",
"10",
"00",
"00",
"01",
"00",
"10",
"10",
"01",
"01",
"10",
"00",
"00",
"00",
"01",
"01",
"01",
"01",
"10",
"01",
"01",
"11",
"11",
"01",
"10",
"00",
"01",
"10",
"00",
"00",
"11",
"00",
"11",
"11",
"01",
"10",
"10",
"01",
"11",
"01",
"10",
"01",
"11",
"11",
"10",
"11",
"01",
"00",
"11",
"11",
"11",
"11",
"01",
"11",
"10",
"10",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"11",
"10",
"01",
"11",
"00",
"10",
"01",
"11",
"01",
"11",
"01",
"11",
"01",
"11",
"10",
"01",
"00",
"00",
"11",
"11",
"00",
"00",
"11",
"00",
"11",
"11",
"11",
"10",
"10",
"10",
"01",
"10",
"11",
"01",
"10",
"01",
"01",
"11",
"00",
"11",
"11",
"11",
"01",
"11",
"11",
"01",
"10",
"11",
"00",
"00",
"00",
"10",
"10",
"10",
"11",
"11",
"01",
"00",
"00",
"00",
"11",
"01",
"10",
"00",
"10",
"11",
"11",
"00",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"00",
"11",
"10",
"00",
"11",
"00",
"00",
"01",
"01",
"00",
"01",
"01",
"10",
"01",
"00",
"10",
"00",
"10",
"11",
"11",
"11",
"01",
"11",
"10",
"01",
"10",
"10",
"00",
"10",
"11",
"01",
"01",
"01",
"11",
"00",
"11",
"00",
"00",
"10",
"11",
"00",
"00",
"00",
"01",
"10",
"10",
"00",
"00",
"11",
"10",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"10",
"00",
"11",
"01",
"01",
"11",
"10",
"01",
"11",
"10",
"01",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"11",
"11",
"00",
"01",
"10",
"11",
"00",
"01",
"00",
"11",
"11",
"11",
"01",
"11",
"00",
"01",
"10",
"00",
"01",
"00",
"10",
"11",
"11",
"10",
"00",
"01",
"11",
"00",
"00",
"00",
"01",
"01",
"00",
"10",
"00",
"11",
"01",
"01",
"00",
"10",
"01",
"11",
"01",
"11",
"01",
"01",
"10",
"11",
"11",
"11",
"00",
"10",
"00",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"00",
"01",
"11",
"11",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"11",
"01",
"11",
"10",
"01",
"01",
"01",
"11",
"10",
"11",
"00",
"00",
"11",
"11",
"11",
"00",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"10",
"01",
"10",
"00",
"00",
"10",
"00",
"11",
"00",
"01",
"00",
"11",
"00",
"01",
"01",
"10",
"11",
"10",
"00",
"11",
"10",
"00",
"11",
"10",
"10",
"10",
"10",
"11",
"01",
"01",
"10",
"01",
"10",
"00",
"01",
"11",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"00",
"11",
"01",
"11",
"10",
"00",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"10",
"00",
"10",
"00",
"11",
"00",
"00",
"11",
"01",
"01",
"10",
"01",
"00",
"11",
"00",
"11",
"01",
"11",
"11",
"00",
"10",
"01",
"00",
"10",
"11",
"01",
"11",
"11",
"10",
"01",
"01",
"00",
"10",
"01",
"11",
"10",
"10",
"10",
"11",
"01",
"11",
"01",
"00",
"00",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"01",
"01",
"01",
"01",
"00",
"10",
"00",
"10",
"01",
"11",
"10",
"01",
"01",
"00",
"01",
"10",
"01",
"10",
"11",
"11",
"11",
"10",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"11",
"00",
"01",
"10",
"11",
"01",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"11",
"00",
"00",
"11",
"00",
"00",
"11",
"11",
"00",
"00",
"11",
"10",
"01",
"11",
"00",
"11",
"10",
"00",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"10",
"00",
"11",
"00",
"01",
"00",
"00",
"10",
"11",
"01",
"10",
"10",
"00",
"01",
"00",
"00",
"11",
"01",
"00",
"00",
"01",
"00",
"11",
"00",
"10",
"00",
"10",
"00",
"11",
"00",
"01",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"00",
"01",
"11",
"11",
"00",
"10",
"11",
"01",
"10",
"01",
"10",
"10",
"00",
"01",
"00",
"11",
"10",
"00",
"11",
"10",
"11",
"11",
"10",
"00",
"11",
"11",
"00",
"10",
"11",
"00",
"10",
"11",
"10",
"11",
"01",
"00",
"00",
"00",
"10",
"00",
"10",
"11",
"00",
"10",
"11",
"10",
"10",
"10",
"10",
"00",
"11",
"01",
"10",
"10",
"11",
"11",
"11",
"00",
"11",
"00",
"11",
"11",
"10",
"01",
"11",
"00",
"01",
"11",
"01",
"01",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"10",
"10",
"10",
"01",
"10",
"00",
"11",
"00",
"10",
"00",
"11",
"00",
"10",
"00",
"10",
"11",
"11",
"10",
"11",
"00",
"10",
"01",
"01",
"11",
"11",
"10",
"10",
"10",
"01",
"01",
"00",
"01",
"11",
"01",
"01",
"10",
"00",
"10",
"11",
"10",
"01",
"11",
"01",
"11",
"01",
"01",
"11",
"01",
"01",
"00",
"11",
"01",
"11",
"00",
"01",
"11",
"11",
"01",
"00",
"01",
"01",
"11",
"00",
"11",
"10",
"01",
"00",
"11",
"01",
"11",
"10",
"01",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"11",
"01",
"10",
"10",
"01",
"11",
"00",
"00",
"01",
"01",
"11",
"10",
"10",
"00",
"10",
"10",
"11",
"10",
"01",
"11",
"00",
"00",
"10",
"00",
"01",
"00",
"01",
"11",
"00",
"11",
"11",
"01",
"11",
"01",
"10",
"10",
"01",
"00",
"10",
"10",
"10",
"00",
"00",
"11",
"00",
"00",
"11",
"10",
"10",
"10",
"10",
"10",
"11",
"10",
"11",
"00",
"01",
"01",
"11",
"01",
"10",
"10",
"01",
"10",
"00",
"10",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"00",
"00",
"01",
"11",
"01",
"01",
"01",
"10",
"10",
"11",
"01",
"01",
"11",
"01",
"11",
"00",
"11",
"10",
"01",
"00",
"11",
"01",
"10",
"11",
"00",
"11",
"10",
"10",
"00",
"01",
"00",
"01",
"10",
"01",
"01",
"11",
"00",
"11",
"01",
"11",
"11",
"10",
"11",
"00",
"10",
"11",
"10",
"11",
"00",
"01",
"10",
"11",
"11",
"10",
"01",
"11",
"01",
"01",
"01",
"11",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"00",
"11",
"10",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"01",
"01",
"00",
"10",
"11",
"11",
"11",
"10",
"00",
"10",
"00",
"11",
"01",
"11",
"00",
"10",
"11",
"00",
"00",
"10",
"01",
"11",
"00",
"11",
"11",
"01",
"10",
"11",
"01",
"10",
"10",
"11",
"01",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"01",
"11",
"00",
"11",
"11",
"01",
"10",
"11",
"11",
"00",
"00",
"01",
"00",
"01",
"10",
"01",
"10",
"00",
"01",
"00",
"01",
"00",
"11",
"11",
"11",
"00",
"00",
"00",
"01",
"00",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"00",
"11",
"01",
"11",
"01",
"10",
"11",
"01",
"10",
"11",
"01",
"11",
"00",
"01",
"00",
"00",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"10",
"01",
"00",
"00",
"10",
"10",
"11",
"00",
"01",
"11",
"01",
"10",
"11",
"00",
"00",
"00",
"10",
"01",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"11",
"00",
"00",
"01",
"11",
"01",
"01",
"01",
"01",
"11",
"11",
"00",
"10",
"01",
"11",
"10",
"00",
"10",
"10",
"10",
"11",
"00",
"01",
"01",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"00",
"11",
"10",
"10",
"01",
"11",
"01",
"11",
"11",
"10",
"00",
"10",
"00",
"11",
"10",
"10",
"01",
"00",
"00",
"01",
"01",
"10",
"11",
"00",
"00",
"10",
"00",
"00",
"01",
"10",
"11",
"01",
"01",
"01",
"10",
"11",
"11",
"01",
"11",
"10",
"00",
"10",
"10",
"00",
"11",
"01",
"00",
"01",
"00",
"00",
"00",
"01",
"11",
"01",
"00",
"01",
"11",
"01",
"11",
"01",
"01",
"00",
"01",
"00",
"11",
"01",
"10",
"11",
"11",
"01",
"00",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"10",
"00",
"10",
"00",
"11",
"11",
"11",
"00",
"00",
"00",
"10",
"00",
"11",
"01",
"00",
"00",
"10",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"00",
"10",
"11",
"11",
"00",
"10",
"01",
"00",
"01",
"11",
"00",
"00",
"01",
"11",
"10",
"10",
"00",
"01",
"11",
"00",
"10",
"00",
"00",
"01",
"11",
"01",
"01",
"11",
"11",
"11",
"10",
"10",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"01",
"01",
"00",
"10",
"00",
"01",
"10",
"10",
"00",
"11",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"10",
"01",
"00",
"11",
"01",
"10",
"10",
"11",
"00",
"00",
"01",
"01",
"00",
"11",
"01",
"11",
"00",
"00",
"11",
"01",
"00",
"01",
"11",
"10",
"01",
"11",
"10",
"01",
"01",
"00",
"01",
"11",
"01",
"11",
"00",
"01",
"00",
"00",
"00",
"01",
"10",
"01",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"00",
"10",
"11",
"01",
"11",
"00",
"11",
"00",
"10",
"00",
"11",
"10",
"10",
"11",
"00",
"01",
"10",
"00",
"00",
"11",
"01",
"10",
"10",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"11",
"01",
"01",
"01",
"00",
"01",
"10",
"10",
"00",
"01",
"00",
"01",
"01",
"01",
"10",
"00",
"00",
"11",
"10",
"11",
"11",
"01",
"00",
"00",
"10",
"10",
"01",
"01",
"01",
"00",
"01",
"10",
"11",
"10",
"01",
"00",
"11",
"01",
"01",
"11",
"01",
"00",
"11",
"10",
"00",
"00",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"01",
"00",
"11",
"01",
"11",
"10",
"00",
"01",
"10",
"01",
"10",
"01",
"10",
"10",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"01",
"00",
"01",
"11",
"00",
"01",
"10",
"00",
"01",
"11",
"00",
"01",
"10",
"00",
"00",
"11",
"10",
"00",
"01",
"00",
"10",
"01",
"10",
"00",
"10",
"10",
"01",
"10",
"10",
"10",
"11",
"10",
"00",
"11",
"10",
"01",
"10",
"10",
"00",
"01",
"10",
"10",
"11",
"11",
"00",
"11",
"11",
"01",
"01",
"00",
"00",
"11",
"10",
"00",
"11",
"01",
"11",
"01",
"11",
"10",
"01",
"01",
"00",
"01",
"11",
"00",
"10",
"10",
"11",
"01",
"00",
"00",
"10",
"11",
"01",
"00",
"10",
"10",
"11",
"11",
"10",
"00",
"01",
"01",
"01",
"00",
"11",
"10",
"01",
"11",
"11",
"10",
"01",
"00",
"11",
"10",
"11",
"00",
"11",
"10",
"10",
"01",
"11",
"10",
"10",
"01",
"11",
"01",
"10",
"10",
"11",
"10",
"00",
"11",
"10",
"10",
"00",
"10",
"11",
"00",
"01",
"00",
"10",
"01",
"00",
"00",
"01",
"11",
"00",
"10",
"00",
"01",
"10",
"00",
"00",
"11",
"10",
"01",
"11",
"10",
"01",
"11",
"10",
"01",
"10",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"11",
"00",
"11",
"10",
"10",
"10",
"01",
"00",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"10",
"11",
"11",
"00",
"11",
"00",
"10",
"01",
"10",
"01",
"11",
"01",
"01",
"10",
"10",
"10",
"10",
"01",
"11",
"01",
"01",
"10",
"01",
"01",
"01",
"11",
"11",
"00",
"11",
"01",
"10",
"11",
"00",
"01",
"01",
"00",
"11",
"01",
"11",
"00",
"10",
"01",
"01",
"00",
"10",
"11",
"01",
"01",
"00",
"11",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"01",
"00",
"01",
"10",
"11",
"11",
"01",
"00",
"11",
"10",
"00",
"01",
"11",
"00",
"11",
"00",
"11",
"01",
"00",
"10",
"11",
"10",
"00",
"00",
"11",
"10",
"10",
"10",
"11",
"11",
"00",
"00",
"10",
"10",
"10",
"00",
"01",
"00",
"10",
"11",
"11",
"11",
"00",
"01",
"11",
"11",
"10",
"10",
"01",
"10",
"00",
"01",
"00",
"11",
"00",
"10",
"11",
"11",
"11",
"11",
"01",
"00",
"11",
"00",
"10",
"00",
"11",
"11",
"11",
"01",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"11",
"01",
"10",
"00",
"00",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"10",
"01",
"10",
"00",
"00",
"11",
"10",
"01",
"10",
"11",
"10",
"10",
"00",
"00",
"01",
"10",
"11",
"00",
"11",
"11",
"11",
"11",
"01",
"00",
"00",
"01",
"11",
"10",
"11",
"11",
"01",
"00",
"10",
"01",
"01",
"11",
"11",
"11",
"00",
"00",
"10",
"01",
"00",
"00",
"00",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"01",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"01",
"00",
"01",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"10",
"00",
"11",
"11",
"11",
"10",
"00",
"10",
"01",
"10",
"11",
"10",
"00",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"11",
"00",
"11",
"01",
"01",
"01",
"01",
"10",
"11",
"10",
"11",
"10",
"01",
"01",
"01",
"10",
"10",
"11",
"10",
"00",
"01",
"10",
"10",
"11",
"11",
"01",
"11",
"11",
"01",
"11",
"00",
"10",
"01",
"01",
"00",
"11",
"11",
"01",
"01",
"11",
"01",
"01",
"00",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"00",
"00",
"01",
"10",
"10",
"11",
"00",
"11",
"11",
"00",
"01",
"11",
"01",
"11",
"01",
"00",
"00",
"00",
"01",
"00",
"10",
"01",
"00",
"11",
"10",
"10",
"11",
"11",
"10",
"00",
"01",
"10",
"00",
"01",
"10",
"01",
"10",
"11",
"01",
"10",
"00",
"01",
"00",
"00",
"11",
"10",
"11",
"10",
"00",
"11",
"00",
"00",
"11",
"11",
"01",
"11",
"10",
"00",
"01",
"00",
"11",
"10",
"10",
"00",
"00",
"01",
"11",
"11",
"01",
"00",
"10",
"01",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"11",
"00",
"00",
"11",
"11",
"00",
"10",
"00",
"10",
"00",
"01",
"01",
"11",
"00",
"00",
"10",
"11",
"01",
"11",
"00",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"00",
"11",
"01",
"00",
"11",
"01",
"00",
"01",
"01",
"00",
"00",
"10",
"00",
"00",
"10",
"10",
"00",
"00",
"10",
"01",
"00",
"10",
"01",
"00",
"01",
"01",
"00",
"00",
"00",
"01",
"11",
"11",
"10",
"11",
"00",
"10",
"01",
"01",
"10",
"11",
"00",
"11",
"11",
"10",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"11",
"00",
"11",
"10",
"01",
"11",
"00",
"10",
"00",
"10",
"01",
"10",
"10",
"00",
"11",
"10",
"11",
"11",
"11",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"00",
"01",
"10",
"01",
"01",
"10",
"10",
"11",
"00",
"00",
"10",
"10",
"01",
"10",
"10",
"11",
"01",
"00",
"11",
"00",
"01",
"11",
"11",
"00",
"00",
"11",
"11",
"11",
"11",
"11",
"01",
"00",
"01",
"01",
"11",
"01",
"10",
"00",
"10",
"00",
"01",
"00",
"00",
"01",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"00",
"10",
"10",
"11",
"10",
"11",
"11",
"10",
"10",
"01",
"00",
"01",
"00",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"00",
"10",
"11",
"01",
"11",
"01",
"00",
"10",
"10",
"11",
"11",
"00",
"00",
"10",
"10",
"11",
"10",
"11",
"01",
"01",
"11",
"11",
"10",
"10",
"01",
"01",
"01",
"00",
"10",
"10",
"00",
"10",
"10",
"00",
"10",
"01",
"11",
"11",
"10",
"00",
"01",
"11",
"11",
"01",
"01",
"01",
"11",
"10",
"01",
"10",
"01",
"10",
"11",
"10",
"11",
"00",
"10",
"00",
"01",
"01",
"10",
"00",
"11",
"00",
"11",
"10",
"10",
"10",
"00",
"10",
"00",
"11",
"11",
"00",
"00",
"10",
"10",
"01",
"10",
"01",
"00",
"10",
"11",
"11",
"00",
"11",
"11",
"10",
"10",
"11",
"01",
"11",
"00",
"01",
"10",
"10",
"10",
"01",
"10",
"00",
"10",
"01",
"00",
"00",
"10",
"10",
"11",
"00",
"10",
"01",
"11",
"01",
"11",
"00",
"11",
"10",
"10",
"01",
"11",
"00",
"01",
"10",
"00",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"00",
"00",
"11",
"00",
"01",
"10",
"10",
"10",
"11",
"11",
"00",
"01",
"11",
"01",
"11",
"10",
"11",
"01",
"01",
"00",
"01",
"00",
"01",
"01",
"00",
"10",
"00",
"10",
"01",
"10",
"00",
"01",
"01",
"00",
"11",
"01",
"11",
"01",
"11",
"11",
"00",
"11",
"01",
"01",
"10",
"10",
"11",
"10",
"00",
"00",
"10",
"01",
"01",
"11",
"11",
"01",
"00",
"00",
"10",
"00",
"00",
"10",
"00",
"10",
"11",
"00",
"11",
"00",
"11",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"11",
"01",
"00",
"00",
"01",
"10",
"10",
"01",
"11",
"00",
"01",
"00",
"01",
"00",
"10",
"01",
"11",
"01",
"01",
"00",
"00",
"01",
"11",
"00",
"01",
"11",
"11",
"00",
"01",
"11",
"10",
"11",
"10",
"11",
"10",
"01",
"10",
"10",
"00",
"00",
"11",
"01",
"00",
"01",
"01",
"11",
"00",
"01",
"00",
"00",
"11",
"11",
"00",
"10",
"10",
"11",
"11",
"01",
"01",
"11",
"01",
"00",
"11",
"01",
"01",
"11",
"10",
"10",
"11",
"01",
"11",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"00",
"10",
"01",
"11",
"00",
"10",
"11",
"10",
"01",
"01",
"10",
"00",
"01",
"01",
"01",
"00",
"01",
"00",
"10",
"01",
"01",
"11",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"11",
"10",
"00",
"01",
"10",
"01",
"00",
"10",
"10",
"01",
"11",
"01",
"00",
"10",
"01",
"10",
"10",
"11",
"01",
"01",
"00",
"10",
"00",
"11",
"11",
"11",
"00",
"10",
"01",
"11",
"10",
"00",
"11",
"00",
"11",
"00",
"11",
"01",
"00",
"10",
"01",
"01",
"11",
"11",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"00",
"11",
"11",
"01",
"11",
"11",
"10",
"01",
"01",
"10",
"00",
"01",
"00",
"10",
"10",
"11",
"11",
"10",
"10",
"00",
"01",
"00",
"11",
"01",
"00",
"11",
"00",
"00",
"00",
"11",
"00",
"01",
"00",
"11",
"11",
"00",
"11",
"11",
"01",
"01",
"10",
"01",
"10",
"01",
"00",
"01",
"11",
"10",
"10",
"00",
"11",
"01",
"01",
"00",
"01",
"01",
"01",
"11",
"00",
"10",
"00",
"01",
"11",
"00",
"00",
"11",
"00",
"10",
"10",
"01",
"10",
"00",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"11",
"00",
"10",
"11",
"01",
"10",
"11",
"11",
"11",
"01",
"11",
"01",
"10",
"01",
"00",
"10",
"10",
"00",
"01",
"11",
"00",
"10",
"11",
"01",
"10",
"11",
"01",
"10",
"11",
"11",
"00",
"10",
"00",
"00",
"01",
"10",
"01",
"00",
"00",
"00",
"11",
"10",
"00",
"11",
"01",
"10",
"01",
"11",
"11",
"01",
"11",
"10",
"11",
"00",
"01",
"11",
"10",
"11",
"00",
"11",
"00",
"11",
"11",
"00",
"11",
"10",
"00",
"10",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"10",
"00",
"01",
"10",
"01",
"01",
"10",
"10",
"01",
"01",
"01",
"00",
"10",
"11",
"01",
"11",
"00",
"01",
"10",
"00",
"10",
"01",
"00",
"10",
"11",
"00",
"01",
"11",
"00",
"01",
"11",
"10",
"11",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"01",
"00",
"01",
"01",
"01",
"01",
"10",
"11",
"00",
"11",
"00",
"11",
"10",
"01",
"00",
"01",
"11",
"10",
"10",
"01",
"01",
"10",
"11",
"00",
"01",
"11",
"01",
"10",
"11",
"01",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"11",
"11",
"01",
"11",
"10",
"01",
"01",
"10",
"11",
"00",
"11",
"10",
"00",
"00",
"10",
"01",
"10",
"11",
"00",
"00",
"11",
"10",
"11",
"11",
"11",
"11",
"11",
"00",
"11",
"01",
"11",
"11",
"10",
"11",
"00",
"00",
"00",
"00",
"11",
"00",
"01",
"11",
"00",
"01",
"10",
"00",
"11",
"11",
"00",
"11",
"10",
"11",
"11",
"11",
"01",
"10",
"11",
"10",
"00",
"00",
"01",
"01",
"11",
"10",
"10",
"00",
"00",
"11",
"11",
"10",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"10",
"01",
"11",
"10",
"11",
"00",
"00",
"11",
"10",
"00",
"00",
"01",
"00",
"00",
"10",
"00",
"11",
"10",
"01",
"00",
"10",
"11",
"10",
"00",
"11",
"01",
"01",
"00",
"01",
"10",
"10",
"11",
"11",
"00",
"00",
"00",
"11",
"10",
"11",
"01",
"10",
"01",
"00",
"00",
"01",
"11",
"01",
"11",
"10",
"00",
"10",
"01",
"11",
"10",
"00",
"00",
"10",
"00",
"01",
"00",
"10",
"00",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"01",
"01",
"00",
"00",
"11",
"11",
"01",
"10",
"11",
"00",
"01",
"10",
"01",
"00",
"01",
"01",
"00",
"01",
"00",
"00",
"00",
"01",
"10",
"10",
"10",
"11",
"11",
"10",
"11",
"10",
"11",
"10",
"00",
"01",
"01",
"11",
"01",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"01",
"01",
"10",
"00",
"01",
"01",
"01",
"10",
"00",
"11",
"11",
"11",
"01",
"11",
"11",
"00",
"01",
"01",
"10",
"00",
"10",
"00",
"11",
"01",
"10",
"01",
"11",
"11",
"01",
"00",
"01",
"01",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"10",
"00",
"01",
"01",
"00",
"10",
"10",
"00",
"00",
"01",
"10",
"01",
"00",
"00",
"00",
"10",
"11",
"00",
"01",
"00",
"01",
"01",
"10",
"10",
"00",
"01",
"10",
"00",
"10",
"10",
"11",
"00",
"00",
"10",
"10",
"10",
"01",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"11",
"00",
"11",
"00",
"11",
"00",
"10",
"00",
"10",
"10",
"10",
"00",
"00",
"11",
"10",
"01",
"00",
"11",
"11",
"10",
"10",
"11",
"11",
"01",
"00",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"00",
"10",
"11",
"00",
"10",
"01",
"00",
"10",
"01",
"10",
"11",
"01",
"11",
"10",
"00",
"01",
"11",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"10",
"10",
"00",
"10",
"10",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"00",
"10",
"00",
"10",
"00",
"11",
"10",
"01",
"10",
"00",
"01",
"10",
"00",
"00",
"01",
"00",
"00",
"11",
"10",
"10",
"11",
"01",
"00",
"00",
"00",
"10",
"00",
"11",
"00",
"11",
"11",
"11",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"00",
"11",
"11",
"11",
"11",
"01",
"10",
"10",
"00",
"01",
"00",
"00",
"10",
"10",
"00",
"10",
"00",
"11",
"11",
"01",
"01",
"10",
"01",
"10",
"00",
"01",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"10",
"00",
"01",
"01",
"01",
"11",
"10",
"11",
"01",
"11",
"01",
"00",
"11",
"01",
"00",
"01",
"10",
"00",
"01",
"10",
"11",
"10",
"00",
"11",
"01",
"10",
"10",
"01",
"01",
"00",
"01",
"01",
"10",
"01",
"01",
"11",
"11",
"01",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"10",
"01",
"00",
"01",
"10",
"01",
"10",
"11",
"00",
"11",
"00",
"11",
"10",
"10",
"11",
"01",
"01",
"10",
"00",
"11",
"01",
"10",
"10",
"10",
"01",
"11",
"00",
"10",
"11",
"11",
"11",
"01",
"00",
"01",
"11",
"10",
"11",
"10",
"10",
"10",
"01",
"00",
"10",
"11",
"00",
"11",
"01",
"01",
"11",
"10",
"00",
"01",
"11",
"10",
"01",
"10",
"10",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"11",
"10",
"01",
"10",
"01",
"01",
"01",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"11",
"10",
"11",
"00",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"11",
"00",
"01",
"01",
"00",
"10",
"00",
"01",
"00",
"11",
"11",
"10",
"00",
"10",
"11",
"11",
"00",
"10",
"10",
"10",
"10",
"01",
"10",
"00",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"00",
"11",
"01",
"01",
"10",
"01",
"00",
"00",
"01",
"01",
"01",
"01",
"10",
"11",
"10",
"10",
"00",
"11",
"01",
"01",
"01",
"10",
"01",
"10",
"10",
"01",
"01",
"00",
"01",
"10",
"01",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"10",
"10",
"01",
"00",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"00",
"01",
"00",
"10",
"01",
"10",
"11",
"00",
"00",
"01",
"11",
"01",
"10",
"01",
"10",
"01",
"00",
"00",
"00",
"11",
"11",
"01",
"01",
"01",
"01",
"10",
"10",
"10",
"11",
"01",
"01",
"10",
"00",
"01",
"00",
"00",
"10",
"00",
"10",
"11",
"10",
"01",
"11",
"10",
"00",
"00",
"10",
"11",
"01",
"00",
"01",
"00",
"10",
"10",
"10",
"11",
"01",
"01",
"00",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"11",
"01",
"00",
"10",
"01",
"11",
"11",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"11",
"00",
"10",
"10",
"10",
"11",
"10",
"01",
"01",
"01",
"11",
"00",
"11",
"00",
"01",
"10",
"11",
"00",
"00",
"11",
"10",
"00",
"00",
"01",
"11",
"10",
"11",
"10",
"01",
"11",
"11",
"00",
"01",
"10",
"10",
"10",
"01",
"00",
"11",
"11",
"00",
"11",
"10",
"11",
"11",
"00",
"00",
"11",
"01",
"11",
"10",
"01",
"10",
"01",
"11",
"01",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"10",
"01",
"01",
"00",
"00",
"11",
"01",
"11",
"01",
"01",
"01",
"00",
"01",
"00",
"10",
"10",
"00",
"11",
"11",
"10",
"11",
"11",
"11",
"01",
"10",
"10",
"11",
"10",
"11",
"10",
"01",
"10",
"10",
"10",
"11",
"10",
"11",
"01",
"01",
"00",
"11",
"01",
"11",
"01",
"00",
"10",
"10",
"10",
"10",
"00",
"10",
"11",
"01",
"01",
"11",
"10",
"00",
"01",
"11",
"01",
"00",
"10",
"01",
"00",
"11",
"01",
"11",
"11",
"00",
"10",
"01",
"01",
"01",
"11",
"00",
"00",
"11",
"01",
"01",
"11",
"01",
"00",
"01",
"01",
"11",
"00",
"01",
"00",
"10",
"10",
"11",
"00",
"11",
"11",
"00",
"01",
"00",
"01",
"00",
"11",
"11",
"00",
"01",
"01",
"00",
"00",
"11",
"10",
"11",
"11",
"00",
"10",
"10",
"11",
"01",
"10",
"11",
"01",
"01",
"01",
"01",
"00",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"01",
"01",
"10",
"11",
"10",
"00",
"11",
"00",
"11",
"10",
"00",
"01",
"10",
"00",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"01",
"11",
"11",
"00",
"11",
"01",
"01",
"10",
"10",
"00",
"11",
"01",
"10",
"01",
"00",
"11",
"11",
"10",
"11",
"11",
"01",
"11",
"10",
"10",
"00",
"01",
"00",
"10",
"01",
"00",
"01",
"00",
"11",
"00",
"11",
"10",
"00",
"10",
"00",
"00",
"01",
"01",
"11",
"00",
"10",
"00",
"11",
"10",
"00",
"10",
"11",
"00",
"11",
"11",
"10",
"00",
"01",
"10",
"01",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"01",
"11",
"00",
"01",
"01",
"01",
"01",
"10",
"00",
"00",
"01",
"10",
"00",
"10",
"10",
"00",
"11",
"10",
"10",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"10",
"11",
"01",
"10",
"00",
"11",
"11",
"10",
"10",
"01",
"01",
"11",
"00",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"01",
"01",
"11",
"00",
"10",
"11",
"01",
"00",
"10",
"10",
"01",
"01",
"01",
"01",
"10",
"01",
"00",
"10",
"10",
"11",
"00",
"10",
"01",
"11",
"10",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"00",
"01",
"00",
"11",
"10",
"00",
"01",
"10",
"00",
"10",
"01",
"00",
"00",
"10",
"00",
"00",
"01",
"11",
"11",
"10",
"00",
"01",
"00",
"00",
"11",
"11",
"10",
"10",
"00",
"00",
"10",
"10",
"10",
"01",
"11",
"01",
"00",
"11",
"00",
"01",
"10",
"01",
"00",
"10",
"00",
"11",
"11",
"00",
"10",
"11",
"01",
"00",
"11",
"11",
"01",
"00",
"01",
"00",
"00",
"00",
"00",
"11",
"00",
"11",
"11",
"10",
"00",
"01",
"00",
"00",
"00",
"01",
"10",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"01",
"00",
"01",
"10",
"01",
"10",
"10",
"00",
"11",
"10",
"00",
"10",
"10",
"10",
"10",
"01",
"10",
"11",
"11",
"01",
"00",
"10",
"00",
"00",
"10",
"10",
"01",
"10",
"00",
"10",
"10",
"11",
"11",
"01",
"00",
"11",
"10",
"11",
"01",
"01",
"10",
"10",
"00",
"10",
"10",
"10",
"01",
"11",
"11",
"10",
"10",
"11",
"11",
"10",
"01",
"11",
"01",
"00",
"00",
"01",
"01",
"01",
"11",
"01",
"00",
"01",
"01",
"10",
"10",
"01",
"00",
"01",
"10",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"10",
"01",
"11",
"11",
"00",
"11",
"01",
"00",
"10",
"00",
"00",
"10",
"00",
"11",
"00",
"10",
"00",
"11",
"10",
"01",
"11",
"00",
"10",
"10",
"11",
"01",
"01",
"11",
"01",
"10",
"01",
"10",
"10",
"10",
"01",
"11",
"01",
"01",
"10",
"00",
"00",
"00",
"01",
"00",
"10",
"11",
"11",
"00",
"00",
"10",
"10",
"01",
"10",
"11",
"10",
"01",
"00",
"11",
"11",
"01",
"00",
"10",
"01",
"00",
"00",
"01",
"11",
"11",
"11",
"01",
"10",
"10",
"11",
"11",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"01",
"00",
"10",
"00",
"00",
"01",
"01",
"11",
"01",
"00",
"10",
"01",
"10",
"11",
"01",
"01",
"11",
"01",
"00",
"10",
"00",
"00",
"00",
"01",
"01",
"00",
"11",
"10",
"01",
"00",
"10",
"11",
"10",
"10",
"00",
"10",
"01",
"11",
"01",
"00",
"11",
"01",
"11",
"01",
"10",
"01",
"01",
"11",
"01",
"11",
"10",
"01",
"01",
"01",
"01",
"11",
"00",
"10",
"11",
"00",
"01",
"11",
"10",
"10",
"11",
"00",
"01",
"11",
"11",
"10",
"01",
"11",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"01",
"10",
"01",
"11",
"00",
"01",
"11",
"10",
"01",
"11",
"00",
"11",
"01",
"10",
"01",
"00",
"11",
"00",
"11",
"00",
"01",
"11",
"10",
"10",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"01",
"10",
"00",
"01",
"01",
"01",
"01",
"00",
"00",
"11",
"00",
"01",
"01",
"10",
"10",
"01",
"00",
"01",
"11",
"01",
"11",
"11",
"01",
"10",
"00",
"00",
"11",
"00",
"00",
"00",
"10",
"01",
"01",
"10",
"10",
"01",
"11",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"00",
"11",
"10",
"00",
"10",
"00",
"11",
"10",
"01",
"01",
"11",
"10",
"10",
"00",
"10",
"11",
"10",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"11",
"11",
"11",
"01",
"10",
"10",
"11",
"11",
"01",
"10",
"00",
"01",
"11",
"10",
"11",
"00",
"10",
"01",
"10",
"00",
"01",
"01",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"00",
"10",
"11",
"11",
"11",
"00",
"10",
"01",
"11",
"00",
"01",
"11",
"00",
"00",
"00",
"10",
"01",
"00",
"00",
"00",
"10",
"01",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"11",
"10",
"00",
"00",
"11",
"00",
"11",
"00",
"00",
"10",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"10",
"11",
"11",
"01",
"11",
"01",
"01",
"00",
"01",
"01",
"11",
"11",
"10",
"10",
"11",
"00",
"11",
"00",
"01",
"11",
"00",
"01",
"01",
"00",
"00",
"11",
"11",
"11",
"11",
"11",
"11",
"11",
"11",
"01",
"10",
"11",
"11",
"11",
"10",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"01",
"10",
"10",
"01",
"01",
"01",
"01",
"00",
"00",
"01",
"01",
"01",
"00",
"00",
"01",
"11",
"00",
"00",
"10",
"01",
"00",
"11",
"11",
"00",
"00",
"01",
"11",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"01",
"10",
"10",
"00",
"01",
"01",
"10",
"00",
"10",
"00",
"00",
"00",
"01",
"01",
"01",
"10",
"01",
"01",
"11",
"00",
"11",
"10",
"00",
"00",
"01",
"10",
"00",
"00",
"10",
"10",
"00",
"00",
"01",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"00",
"00",
"00",
"00",
"11",
"00",
"11",
"00",
"00",
"00",
"11",
"10",
"00",
"11",
"00",
"11",
"01",
"11",
"10",
"10",
"10",
"11",
"11",
"11",
"01",
"10",
"00",
"10",
"00",
"00",
"01",
"10",
"01",
"10",
"10",
"10",
"11",
"00",
"11",
"01",
"01",
"00",
"01",
"10",
"00",
"00",
"10",
"11",
"01",
"10",
"11",
"01",
"01",
"11",
"00",
"01",
"01",
"10",
"00",
"01",
"11",
"11",
"00",
"11",
"00",
"10",
"11",
"00",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"10",
"10",
"10",
"11",
"11",
"10",
"00",
"00",
"01",
"01",
"00",
"01",
"11",
"10",
"00",
"10",
"11",
"10",
"10",
"01",
"11",
"11",
"11",
"00",
"01",
"00",
"00",
"10",
"10",
"01",
"11",
"00",
"10",
"00",
"11",
"00",
"11",
"01",
"11",
"11",
"10",
"10",
"00",
"01",
"00",
"00",
"11",
"11",
"10",
"11",
"00",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"10",
"01",
"10",
"10",
"01",
"10",
"00",
"11",
"01",
"00",
"01",
"00",
"10",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"10",
"00",
"00",
"10",
"01",
"01",
"01",
"00",
"11",
"00",
"01",
"01",
"11",
"10",
"00",
"10",
"11",
"10",
"00",
"11",
"01",
"01",
"00",
"00",
"01",
"11",
"00",
"00",
"11",
"01",
"01",
"01",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"11",
"00",
"10",
"00",
"10",
"01",
"00",
"10",
"10",
"10",
"00",
"10",
"11",
"00",
"11",
"11",
"01",
"10",
"01",
"11",
"00",
"10",
"11",
"00",
"00",
"00",
"11",
"11",
"01",
"00",
"01",
"10",
"11",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"11",
"00",
"10",
"11",
"00",
"10",
"11",
"00",
"00",
"10",
"11",
"00",
"10",
"10",
"00",
"01",
"00",
"10",
"10",
"10",
"01",
"01",
"10",
"00",
"01",
"10",
"01",
"11",
"01",
"00",
"11",
"00",
"01",
"10",
"10",
"10",
"01",
"01",
"01",
"10",
"00",
"10",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"10",
"10",
"10",
"01",
"01",
"11",
"01",
"00",
"01",
"11",
"11",
"10",
"00",
"00",
"10",
"00",
"11",
"11",
"10",
"01",
"01",
"10",
"00",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"11",
"10",
"00",
"11",
"00",
"01",
"00",
"11",
"11",
"01",
"01",
"00",
"00",
"00",
"10",
"00",
"00",
"00",
"10",
"00",
"01",
"01",
"10",
"11",
"11",
"11",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"10",
"00",
"11",
"00",
"01",
"01",
"11",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"00",
"00",
"11",
"10",
"11",
"01",
"01",
"11",
"00",
"11",
"11",
"00",
"11",
"10",
"00",
"11",
"10",
"10",
"10",
"11",
"00",
"00",
"11",
"01",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"00",
"01",
"11",
"01",
"00",
"10",
"10",
"01",
"10",
"00",
"01",
"01",
"00",
"00",
"00",
"11",
"00",
"11",
"01",
"10",
"11",
"00",
"11",
"01",
"01",
"10",
"00",
"11",
"10",
"00",
"10",
"11",
"11",
"00",
"11",
"10",
"00",
"10",
"10",
"10",
"11",
"00",
"01",
"01",
"01",
"10",
"11",
"10",
"01",
"10",
"01",
"01",
"11",
"11",
"10",
"01",
"10",
"10",
"00",
"00",
"01",
"01",
"10",
"11",
"11",
"11",
"10",
"00",
"01",
"00",
"00",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"11",
"10",
"00",
"01",
"11",
"10",
"11",
"01",
"11",
"10",
"00",
"01",
"00",
"01",
"00",
"10",
"10",
"10",
"01",
"10",
"11",
"11",
"11",
"10",
"01",
"11",
"01",
"01",
"00",
"11",
"10",
"00",
"10",
"10",
"01",
"01",
"01",
"01",
"00",
"00",
"01",
"11",
"00",
"00",
"10",
"10",
"01",
"11",
"11",
"11",
"00",
"10",
"10",
"10",
"00",
"11",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"10",
"10",
"10",
"00",
"00",
"00",
"10",
"00",
"00",
"00",
"11",
"01",
"01",
"00",
"11",
"11",
"00",
"00",
"01",
"10",
"10",
"01",
"00",
"00",
"10",
"10",
"00",
"11",
"10",
"01",
"10",
"10",
"01",
"10",
"11",
"10",
"00",
"01",
"01",
"00",
"11",
"11",
"01",
"00",
"01",
"11",
"10",
"11",
"10",
"10",
"00",
"11",
"10",
"01",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"11",
"10",
"00",
"11",
"10",
"01",
"01",
"10",
"11",
"01",
"10",
"01",
"01",
"10",
"01",
"11",
"11",
"11",
"11",
"00",
"00",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"11",
"11",
"00",
"01",
"00",
"11",
"01",
"01",
"00",
"10",
"00",
"10",
"01",
"11",
"01",
"11",
"01",
"01",
"00",
"00",
"00",
"10",
"10",
"01",
"00",
"00",
"11",
"10",
"01",
"11",
"11",
"01",
"11",
"10",
"00",
"10",
"00",
"01",
"11",
"11",
"00",
"01",
"00",
"01",
"11",
"10",
"01",
"11",
"11",
"00",
"00",
"01",
"01",
"00",
"10",
"11",
"00",
"11",
"11",
"10",
"01",
"01",
"01",
"10",
"10",
"00",
"10",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"00",
"00",
"01",
"00",
"01",
"10",
"00",
"10",
"10",
"01",
"01",
"10",
"11",
"00",
"11",
"00",
"00",
"10",
"10",
"11",
"11",
"11",
"01",
"01",
"11",
"01",
"11",
"11",
"00",
"00",
"00",
"01",
"01",
"00",
"00",
"00",
"10",
"00",
"00",
"01",
"01",
"10",
"11",
"00",
"01",
"01",
"00",
"11",
"00",
"00",
"01",
"10",
"01",
"10",
"01",
"10",
"11",
"01",
"01",
"11",
"11",
"11",
"10",
"10",
"01",
"11",
"00",
"11",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"11",
"01",
"10",
"11",
"01",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"01",
"01",
"10",
"00",
"10",
"11",
"00",
"10",
"11",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"00",
"10",
"10",
"11",
"00",
"10",
"00",
"11",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"00",
"00",
"00",
"10",
"00",
"01",
"11",
"00",
"00",
"01",
"11",
"00",
"00",
"01",
"00",
"10",
"00",
"00",
"10",
"01",
"11",
"00",
"10",
"11",
"00",
"00",
"11",
"11",
"10",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"01",
"10",
"10",
"00",
"01",
"01",
"00",
"11",
"01",
"10",
"01",
"01",
"11",
"11",
"11",
"10",
"01",
"00",
"11",
"10",
"01",
"10",
"10",
"10",
"01",
"10",
"01",
"00",
"00",
"00",
"11",
"01",
"00",
"10",
"00",
"00",
"11",
"11",
"00",
"10",
"11",
"00",
"11",
"11",
"01",
"01",
"11",
"01",
"00",
"00",
"01",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"00",
"01",
"01",
"10",
"10",
"00",
"01",
"10",
"01",
"00",
"11",
"01",
"11",
"01",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"10",
"10",
"01",
"11",
"11",
"11",
"00",
"01",
"00",
"00",
"10",
"01",
"11",
"10",
"11",
"11",
"11",
"11",
"11",
"10",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"10",
"01",
"11",
"01",
"01",
"00",
"01",
"11",
"11",
"11",
"00",
"10",
"10",
"11",
"11",
"00",
"11",
"11",
"10",
"10",
"00",
"00",
"01",
"01",
"00",
"01",
"11",
"11",
"00",
"11",
"10",
"01",
"11",
"00",
"01",
"10",
"10",
"00",
"01",
"10",
"01",
"10",
"01",
"10",
"00",
"11",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"00",
"11",
"11",
"10",
"11",
"11",
"01",
"01",
"00",
"11",
"00",
"01",
"11",
"11",
"01",
"10",
"01",
"10",
"00",
"00",
"11",
"01",
"11",
"10",
"10",
"10",
"00",
"10",
"00",
"10",
"10",
"01",
"01",
"00",
"00",
"01",
"01",
"10",
"00",
"01",
"01",
"01",
"10",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"01",
"00",
"10",
"11",
"00",
"10",
"11",
"11",
"01",
"00",
"10",
"01",
"11",
"01",
"10",
"11",
"10",
"10",
"11",
"10",
"11",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"11",
"11",
"01",
"01",
"00",
"11",
"11",
"01",
"00",
"10",
"11",
"10",
"00",
"11",
"11",
"01",
"01",
"11",
"11",
"10",
"11",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"11",
"00",
"10",
"00",
"00",
"01",
"01",
"00",
"01",
"11",
"11",
"10",
"01",
"10",
"01",
"00",
"11",
"00",
"11",
"01",
"11",
"11",
"11",
"00",
"00",
"01",
"10",
"11",
"10",
"10",
"11",
"01",
"10",
"10",
"10",
"10",
"01",
"00",
"10",
"11",
"00",
"10",
"10",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"01",
"00",
"01",
"10",
"01",
"10",
"11",
"00",
"11",
"10",
"01",
"00",
"10",
"01",
"00",
"11",
"01",
"11",
"10",
"11",
"11",
"00",
"11",
"00",
"01",
"01",
"10",
"01",
"11",
"10",
"00",
"11",
"10",
"11",
"00",
"11",
"10",
"00",
"10",
"10",
"01",
"11",
"11",
"10",
"00",
"00",
"01",
"11",
"11",
"01",
"00",
"11",
"00",
"00",
"01",
"11",
"10",
"01",
"11",
"00",
"11",
"10",
"11",
"00",
"00",
"00",
"11",
"00",
"01",
"00",
"01",
"01",
"01",
"11",
"11",
"10",
"11",
"00",
"00",
"00",
"01",
"11",
"11",
"01",
"00",
"10",
"00",
"11",
"01",
"10",
"10",
"01",
"10",
"00",
"01",
"11",
"01",
"11",
"10",
"00",
"01",
"10",
"10",
"10",
"01",
"10",
"10",
"01",
"00",
"10",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"11",
"00",
"01",
"10",
"11",
"00",
"00",
"01",
"10",
"01",
"00",
"11",
"00",
"00",
"11",
"10",
"00",
"01",
"10",
"11",
"11",
"00",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"00",
"00",
"11",
"00",
"11",
"00",
"11",
"01",
"11",
"00",
"01",
"11",
"00",
"10",
"01",
"11",
"00",
"00",
"01",
"00",
"10",
"10",
"00",
"01",
"11",
"01",
"11",
"11",
"10",
"10",
"00",
"00",
"10",
"10",
"00",
"01",
"01",
"10",
"00",
"00",
"00",
"01",
"00",
"00",
"10",
"01",
"00",
"10",
"11",
"10",
"01",
"00",
"01",
"11",
"11",
"10",
"11",
"10",
"00",
"00",
"11",
"10",
"11",
"01",
"11",
"00",
"10",
"00",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"01",
"00",
"00",
"00",
"11",
"00",
"00",
"00",
"11",
"11",
"01",
"01",
"01",
"11",
"00",
"10",
"11",
"11",
"10",
"10",
"01",
"10",
"11",
"10",
"01",
"00",
"11",
"01",
"11",
"11",
"10",
"01",
"10",
"10",
"10",
"01",
"11",
"00",
"01",
"10",
"00",
"11",
"00",
"01",
"11",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"00",
"11",
"00",
"01",
"10",
"10",
"11",
"00",
"11",
"01",
"00",
"01",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"01",
"00",
"11",
"00",
"01",
"01",
"10",
"01",
"11",
"00",
"01",
"10",
"10",
"10",
"00",
"00",
"10",
"00",
"01",
"11",
"11",
"01",
"01",
"00",
"00",
"00",
"10",
"11",
"11",
"10",
"11",
"01",
"00",
"11",
"10",
"00",
"10",
"00",
"10",
"11",
"10",
"00",
"11",
"10",
"11",
"11",
"01",
"11",
"11",
"10",
"00",
"10",
"10",
"00",
"00",
"00",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"10",
"01",
"11",
"00",
"11",
"10",
"11",
"11",
"00",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"00",
"00",
"00",
"00",
"01",
"10",
"11",
"11",
"00",
"10",
"00",
"10",
"00",
"10",
"10",
"10",
"01",
"10",
"11",
"11",
"10",
"11",
"11",
"10",
"01",
"00",
"01",
"00",
"00",
"11",
"10",
"11",
"10",
"11",
"11",
"10",
"10",
"11",
"01",
"01",
"00",
"00",
"01",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"01",
"11",
"11",
"01",
"00",
"10",
"01",
"00",
"10",
"11",
"00",
"01",
"11",
"00",
"00",
"10",
"11",
"01",
"10",
"00",
"11",
"00",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"00",
"01",
"10",
"01",
"00",
"01",
"00",
"10",
"11",
"11",
"11",
"10",
"01",
"11",
"10",
"00",
"10",
"10",
"00",
"00",
"00",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"01",
"11",
"01",
"01",
"10",
"11",
"11",
"11",
"10",
"10",
"01",
"01",
"01",
"00",
"00",
"01",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"11",
"10",
"11",
"01",
"01",
"00",
"11",
"01",
"10",
"11",
"10",
"00",
"01",
"10",
"10",
"10",
"11",
"00",
"01",
"11",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"00",
"10",
"00",
"00",
"00",
"11",
"00",
"00",
"11",
"00",
"11",
"00",
"00",
"11",
"10",
"01",
"01",
"11",
"00",
"00",
"11",
"11",
"11",
"10",
"11",
"00",
"01",
"00",
"11",
"01",
"10",
"01",
"10",
"11",
"10",
"11",
"10",
"11",
"00",
"01",
"00",
"00",
"00",
"10",
"00",
"11",
"11",
"01",
"00",
"01",
"10",
"00",
"11",
"11",
"00",
"00",
"00",
"00",
"01",
"00",
"10",
"01",
"10",
"10",
"00",
"01",
"00",
"00",
"00",
"00",
"11",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"11",
"10",
"00",
"11",
"01",
"01",
"10",
"01",
"01",
"10",
"00",
"01",
"10",
"10",
"10",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"01",
"00",
"00",
"00",
"11",
"10",
"00",
"10",
"01",
"10",
"01",
"00",
"00",
"10",
"00",
"11",
"11",
"01",
"00",
"01",
"01",
"00",
"10",
"10",
"11",
"10",
"11",
"00",
"00",
"11",
"11",
"01",
"00",
"01",
"00",
"01",
"00",
"00",
"00",
"01",
"11",
"11",
"01",
"10",
"10",
"10",
"10",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"10",
"01",
"11",
"00",
"01",
"01",
"00",
"00",
"10",
"01",
"11",
"10",
"10",
"01",
"00",
"11",
"10",
"00",
"11",
"11",
"10",
"11",
"00",
"10",
"00",
"00",
"10",
"11",
"11",
"01",
"01",
"11",
"01",
"10",
"10",
"00",
"00",
"10",
"01",
"11",
"11",
"10",
"11",
"00",
"10",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"11",
"11",
"11",
"10",
"10",
"00",
"10",
"01",
"01",
"01",
"11",
"01",
"10",
"01",
"10",
"01",
"11",
"11",
"10",
"10",
"01",
"01",
"11",
"10",
"10",
"00",
"10",
"00",
"01",
"00",
"11",
"11",
"00",
"11",
"00",
"00",
"01",
"01",
"00",
"11",
"01",
"10",
"11",
"00",
"01",
"00",
"11",
"01",
"10",
"01",
"00",
"10",
"10",
"11",
"11",
"01",
"01",
"00",
"11",
"11",
"11",
"01",
"01",
"11",
"11",
"10",
"01",
"01",
"11",
"00",
"00",
"11",
"10",
"01",
"10",
"00",
"00",
"11",
"10",
"01",
"00",
"01",
"00",
"11",
"11",
"11",
"01",
"01",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"11",
"10",
"11",
"10",
"01",
"10",
"11",
"11",
"00",
"10",
"01",
"00",
"10",
"00",
"10",
"01",
"01",
"11",
"11",
"11",
"11",
"11",
"01",
"10",
"00",
"00",
"10",
"10",
"00",
"00",
"10",
"10",
"11",
"01",
"01",
"11",
"10",
"00",
"01",
"11",
"00",
"01",
"00",
"00",
"10",
"00",
"10",
"11",
"10",
"11",
"01",
"00",
"00",
"10",
"00",
"10",
"00",
"01",
"01",
"01",
"00",
"10",
"01",
"10",
"11",
"00",
"10",
"11",
"01",
"11",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"01",
"00",
"10",
"00",
"11",
"10",
"01",
"11",
"10",
"10",
"11",
"11",
"10",
"00",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"00",
"11",
"01",
"01",
"01",
"10",
"10",
"00",
"00",
"01",
"00",
"10",
"11",
"00",
"10",
"01",
"11",
"00",
"11",
"10",
"00",
"00",
"01",
"11",
"10",
"10",
"01",
"00",
"01",
"01",
"10",
"00",
"11",
"10",
"00",
"11",
"11",
"10",
"10",
"10",
"01",
"10",
"00",
"00",
"10",
"01",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"00",
"00",
"00",
"01",
"11",
"10",
"00",
"11",
"10",
"01",
"11",
"11",
"10",
"00",
"00",
"00",
"00",
"11",
"00",
"11",
"01",
"01",
"10",
"01",
"01",
"00",
"00",
"00",
"01",
"00",
"10",
"10",
"00",
"00",
"01",
"00",
"11",
"00",
"10",
"00",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"00",
"11",
"10",
"10",
"00",
"10",
"00",
"11",
"00",
"01",
"10",
"01",
"10",
"00",
"10",
"01",
"01",
"01",
"01",
"10",
"11",
"01",
"01",
"00",
"00",
"10",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"11",
"10",
"10",
"00",
"00",
"10",
"11",
"11",
"11",
"11",
"00",
"00",
"10",
"10",
"01",
"00",
"11",
"00",
"00",
"11",
"01",
"11",
"11",
"10",
"11",
"11",
"00",
"10",
"01",
"00",
"01",
"11",
"10",
"10",
"00",
"10",
"11",
"00",
"11",
"01",
"10",
"11",
"10",
"00",
"01",
"00",
"00",
"01",
"00",
"10",
"01",
"10",
"11",
"00",
"11",
"11",
"11",
"01",
"10",
"11",
"11",
"10",
"10",
"00",
"11",
"00",
"01",
"10",
"01",
"11",
"10",
"11",
"01",
"11",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"11",
"01",
"00",
"11",
"01",
"00",
"00",
"10",
"00",
"01",
"00",
"01",
"00",
"10",
"01",
"00",
"11",
"00",
"01",
"11",
"00",
"11",
"00",
"01",
"00",
"10",
"00",
"00",
"01",
"00",
"11",
"11",
"11",
"10",
"01",
"00",
"00",
"11",
"01",
"10",
"11",
"00",
"00",
"00",
"10",
"10",
"11",
"00",
"11",
"10",
"11",
"11",
"00",
"01",
"11",
"00",
"00",
"01",
"11",
"10",
"00",
"11",
"00",
"10",
"10",
"10",
"10",
"01",
"01",
"00",
"11",
"01",
"01",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"11",
"01",
"11",
"10",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"00",
"10",
"01",
"10",
"00",
"11",
"01",
"10",
"01",
"00",
"11",
"00",
"10",
"00",
"11",
"00",
"10",
"11",
"10",
"11",
"11",
"01",
"01",
"10",
"10",
"11",
"00",
"00",
"11",
"10",
"01",
"01",
"01",
"11",
"01",
"00",
"01",
"01",
"10",
"00",
"00",
"10",
"01",
"01",
"10",
"00",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"00",
"00",
"00",
"11",
"00",
"01",
"10",
"00",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"01",
"00",
"10",
"00",
"11",
"11",
"00",
"10",
"10",
"00",
"01",
"11",
"01",
"11",
"01",
"00",
"00",
"11",
"11",
"01",
"10",
"11",
"11",
"11",
"01",
"10",
"01",
"10",
"01",
"00",
"11",
"01",
"01",
"00",
"01",
"00",
"00",
"00",
"00",
"01",
"00",
"10",
"10",
"00",
"00",
"10",
"10",
"11",
"11",
"10",
"11",
"10",
"11",
"11",
"10",
"11",
"11",
"01",
"00",
"00",
"00",
"00",
"01",
"01",
"00",
"10",
"11",
"00",
"00",
"01",
"01",
"11",
"01",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"10",
"10",
"11",
"10",
"00",
"10",
"10",
"01",
"00",
"11",
"10",
"11",
"11",
"10",
"11",
"00",
"00",
"10",
"01",
"10",
"10",
"10",
"00",
"10",
"10",
"11",
"11",
"10",
"11",
"00",
"01",
"11",
"00",
"11",
"11",
"00",
"11",
"11",
"01",
"01",
"00",
"00",
"10",
"01",
"10",
"01",
"00",
"11",
"01",
"11",
"00",
"01",
"01",
"00",
"10",
"01",
"10",
"11",
"01",
"01",
"10",
"01",
"10",
"00",
"01",
"11",
"11",
"01",
"10",
"10",
"10",
"10",
"10",
"11",
"11",
"01",
"00",
"00",
"10",
"10",
"01",
"01",
"10",
"10",
"11",
"10",
"01",
"10",
"11",
"01",
"01",
"01",
"11",
"10",
"00",
"10",
"01",
"10",
"11",
"00",
"11",
"00",
"11",
"00",
"00",
"00",
"00",
"01",
"00",
"00",
"01",
"11",
"00",
"00",
"11",
"01",
"10",
"10",
"01",
"10",
"01",
"00",
"01",
"11",
"00",
"11",
"00",
"11",
"00",
"10",
"01",
"10",
"01",
"11",
"10",
"10",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"00",
"11",
"11",
"11",
"10",
"00",
"00",
"01",
"00",
"11",
"00",
"10",
"10",
"10",
"00",
"01",
"00",
"10",
"00",
"01",
"11",
"00",
"11",
"10",
"11",
"10",
"00",
"11",
"00",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"00",
"10",
"10",
"11",
"00",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"01",
"01",
"10",
"00",
"11",
"01",
"10",
"00",
"11",
"00",
"10",
"00",
"00",
"11",
"01",
"00",
"10",
"11",
"11",
"11",
"11",
"10",
"00",
"00",
"10",
"10",
"01",
"00",
"00",
"10",
"01",
"00",
"01",
"01",
"00",
"11",
"01",
"10",
"01",
"01",
"00",
"00",
"00",
"10",
"00",
"10",
"01",
"10",
"00",
"00",
"10",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"10",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"01",
"01",
"00",
"10",
"10",
"01",
"01",
"01",
"10",
"01",
"01",
"00",
"00",
"01",
"11",
"00",
"01",
"10",
"11",
"00",
"11",
"11",
"01",
"10",
"01",
"01",
"10",
"00",
"11",
"00",
"11",
"11",
"10",
"00",
"00",
"00",
"01",
"00",
"00",
"10",
"01",
"10",
"10",
"11",
"01",
"10",
"11",
"11",
"01",
"00",
"00",
"10",
"11",
"10",
"11",
"01",
"01",
"00",
"01",
"10",
"01",
"00",
"01",
"11",
"11",
"10",
"10",
"01",
"10",
"00",
"11",
"10",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"11",
"10",
"10",
"11",
"10",
"00",
"01",
"11",
"11",
"00",
"00",
"00",
"01",
"00",
"00",
"11",
"11",
"10",
"00",
"00",
"01",
"00",
"00",
"01",
"11",
"01",
"00",
"00",
"11",
"10",
"01",
"00",
"00",
"11",
"11",
"11",
"10",
"10",
"00",
"00",
"11",
"00",
"11",
"00",
"00",
"00",
"11",
"00",
"01",
"10",
"00",
"00",
"11",
"10",
"10",
"00",
"00",
"11",
"10",
"00",
"11",
"01",
"10",
"01",
"01",
"00",
"01",
"00",
"00",
"10",
"00",
"01",
"10",
"00",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"10",
"10",
"10",
"10",
"10",
"01",
"01",
"00",
"01",
"11",
"01",
"00",
"01",
"00",
"10",
"11",
"10",
"11",
"00",
"11",
"01",
"01",
"11",
"10",
"01",
"01",
"00",
"01",
"00",
"00",
"10",
"11",
"10",
"00",
"00",
"01",
"10",
"01",
"01",
"00",
"00",
"11",
"10",
"00",
"01",
"00",
"11",
"10",
"10",
"00",
"00",
"10",
"11",
"10",
"01",
"11",
"10",
"01",
"00",
"10",
"00",
"01",
"10",
"00",
"00",
"11",
"10",
"10",
"10",
"00",
"00",
"10",
"11",
"10",
"10",
"11",
"10",
"10",
"00",
"10",
"11",
"01",
"00",
"10",
"00",
"10",
"11",
"01",
"10",
"01",
"00",
"10",
"01",
"10",
"00",
"00",
"01",
"00",
"11",
"01",
"00",
"01",
"10",
"00",
"00",
"11",
"01",
"00",
"00",
"10",
"11",
"11",
"00",
"00",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"00",
"01",
"00",
"11",
"01",
"10",
"01",
"10",
"01",
"10",
"10",
"10",
"10",
"10",
"00",
"00",
"01",
"01",
"10",
"00",
"01",
"10",
"10",
"11",
"00",
"01",
"11",
"01",
"11",
"00",
"11",
"01",
"10",
"01",
"10",
"01",
"10",
"01",
"00",
"11",
"00",
"01",
"00",
"11",
"10",
"01",
"10",
"01",
"10",
"10",
"10",
"00",
"11",
"11",
"01",
"00",
"11",
"11",
"00",
"01",
"11",
"11",
"11",
"01",
"01",
"10",
"00",
"11",
"11",
"11",
"11",
"00",
"10",
"00",
"10",
"00",
"10",
"01",
"00",
"00",
"00",
"10",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"11",
"11",
"10",
"01",
"00",
"00",
"10",
"01",
"11",
"11",
"11",
"01",
"01",
"00",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"11",
"01",
"11",
"01",
"11",
"00",
"00",
"00",
"11",
"11",
"01",
"00",
"01",
"10",
"01",
"00",
"11",
"10",
"01",
"00",
"01",
"00",
"10",
"00",
"11",
"01",
"00",
"00",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"11",
"00",
"11",
"11",
"10",
"01",
"00",
"01",
"01",
"10",
"11",
"11",
"01",
"10",
"00",
"01",
"10",
"11",
"01",
"10",
"10",
"11",
"01",
"11",
"10",
"10",
"00",
"00",
"10",
"01",
"01",
"10",
"01",
"10",
"11",
"10",
"11",
"00",
"00",
"00",
"00",
"10",
"10",
"00",
"11",
"01",
"01",
"11",
"11",
"00",
"10",
"11",
"01",
"01",
"00",
"11",
"11",
"00",
"11",
"10",
"00",
"01",
"10",
"01",
"11",
"00",
"10",
"11",
"00",
"11",
"11",
"00",
"00",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"01",
"01",
"01",
"01",
"01",
"00",
"01",
"11",
"10",
"11",
"11",
"00",
"10",
"11",
"00",
"01",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"00",
"11",
"01",
"11",
"00",
"00",
"11",
"11",
"11",
"10",
"00",
"11",
"00",
"10",
"11",
"10",
"11",
"01",
"00",
"01",
"10",
"00",
"10",
"10",
"00",
"00",
"11",
"11",
"00",
"10",
"01",
"10",
"10",
"00",
"00",
"00",
"10",
"00",
"00",
"10",
"10",
"10",
"10",
"11",
"01",
"11",
"10",
"00",
"10",
"11",
"11",
"11",
"01",
"11",
"00",
"00",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"11",
"00",
"11",
"01",
"00",
"11",
"11",
"10",
"01",
"01",
"11",
"11",
"01",
"10",
"10",
"00",
"00",
"01",
"11",
"10",
"00",
"00",
"10",
"11",
"00",
"11",
"00",
"10",
"11",
"10",
"01",
"00",
"11",
"11",
"00",
"11",
"10",
"10",
"01",
"10",
"00",
"10",
"00",
"01",
"00",
"10",
"11",
"00",
"11",
"11",
"00",
"10",
"01",
"10",
"00",
"00",
"01",
"00",
"10",
"01",
"01",
"01",
"00",
"01",
"00",
"00",
"00",
"11",
"10",
"11",
"10",
"00",
"01",
"10",
"00",
"01",
"01",
"01",
"01",
"11",
"01",
"10",
"11",
"10",
"11",
"11",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"10",
"10",
"01",
"01",
"00",
"11",
"11",
"10",
"11",
"10",
"00",
"10",
"11",
"00",
"00",
"01",
"01",
"10",
"01",
"01",
"01",
"00",
"10",
"01",
"00",
"00",
"00",
"00",
"01",
"10",
"11",
"01",
"01",
"11",
"10",
"01",
"10",
"00",
"01",
"01",
"00",
"01",
"10",
"01",
"00",
"00",
"01",
"01",
"11",
"11",
"10",
"01",
"01",
"00",
"00",
"11",
"00",
"00",
"01",
"01",
"00",
"00",
"00",
"10",
"01",
"10",
"10",
"00",
"11",
"11",
"00",
"00",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"11",
"01",
"11",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"10",
"10",
"10",
"10",
"00",
"11",
"11",
"10",
"10",
"01",
"00",
"00",
"00",
"01",
"10",
"10",
"00",
"10",
"10",
"11",
"00",
"01",
"00",
"00",
"11",
"11",
"11",
"01",
"11",
"00",
"00",
"00",
"11",
"10",
"01",
"00",
"01",
"01",
"00",
"10",
"01",
"11",
"00",
"10",
"01",
"11",
"10",
"11",
"01",
"00",
"01",
"00",
"00",
"01",
"00",
"10",
"10",
"01",
"00",
"11",
"00",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"11",
"00",
"10",
"10",
"11",
"11",
"11",
"01",
"01",
"10",
"11",
"01",
"01",
"01",
"11",
"01",
"10",
"10",
"00",
"10",
"01",
"11",
"00",
"01",
"01",
"11",
"00",
"11",
"11",
"01",
"00",
"10",
"10",
"10",
"10",
"11",
"11",
"10",
"00",
"00",
"01",
"01",
"11",
"00",
"00",
"10",
"10",
"10",
"11",
"00",
"10",
"10",
"10",
"11",
"00",
"00",
"00",
"10",
"01",
"01",
"00",
"11",
"10",
"01",
"11",
"11",
"10",
"00",
"01",
"11",
"00",
"11",
"00",
"10",
"01",
"10",
"10",
"10",
"10",
"01",
"10",
"11",
"00",
"10",
"00",
"00",
"00",
"10",
"11",
"01",
"00",
"00",
"11",
"11",
"11",
"00",
"00",
"10",
"10",
"10",
"00",
"01",
"00",
"10",
"01",
"01",
"11",
"00",
"11",
"11",
"10",
"01",
"00",
"00",
"00",
"10",
"11",
"01",
"10",
"00",
"10",
"11",
"00",
"01",
"01",
"01",
"00",
"10",
"11",
"00",
"11",
"00",
"01",
"01",
"10",
"11",
"10",
"01",
"00",
"01",
"10",
"00",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"10",
"11",
"01",
"01",
"10",
"11",
"00",
"01",
"00",
"10",
"00",
"00",
"00",
"10",
"10",
"01",
"00",
"00",
"10",
"11",
"11",
"01",
"00",
"00",
"11",
"01",
"01",
"10",
"00",
"01",
"10",
"00",
"01",
"00",
"01",
"11",
"11",
"11",
"10",
"11",
"00",
"11",
"01",
"11",
"01",
"11",
"10",
"00",
"00",
"11",
"10",
"11",
"01",
"11",
"01",
"10",
"01",
"00",
"11",
"00",
"00",
"00",
"10",
"11",
"01",
"01",
"00",
"10",
"10",
"00",
"11",
"01",
"10",
"00",
"11",
"11",
"10",
"10",
"11",
"00",
"00",
"01",
"00",
"00",
"00",
"11",
"10",
"00",
"01",
"01",
"10",
"01",
"10",
"11",
"01",
"11",
"10",
"01",
"01",
"01",
"10",
"11",
"00",
"10",
"00",
"01",
"00",
"11",
"10",
"01",
"10",
"00",
"10",
"11",
"01",
"11",
"10",
"10",
"10",
"11",
"00",
"01",
"00",
"01",
"00",
"01",
"01",
"01",
"00",
"10",
"10",
"01",
"00",
"01",
"00",
"01",
"10",
"11",
"11",
"11",
"11",
"01",
"11",
"11",
"00",
"10",
"01",
"10",
"00",
"00",
"00",
"00",
"10",
"00",
"11",
"11",
"00",
"11",
"01",
"01",
"11",
"00",
"01",
"00",
"01",
"11",
"00",
"10",
"10",
"11",
"10",
"00",
"10",
"00",
"10",
"11",
"10",
"01",
"00",
"11",
"10",
"01",
"11",
"10",
"11",
"00",
"11",
"10",
"10",
"01",
"11",
"10",
"00",
"11",
"11",
"10",
"01",
"01",
"00",
"10",
"01",
"11",
"01",
"01",
"01",
"00",
"11",
"01",
"01",
"01",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"10",
"11",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"01",
"10",
"10",
"00",
"11",
"10",
"00",
"00",
"00",
"00",
"10",
"01",
"01",
"00",
"11",
"01",
"00",
"01",
"00",
"11",
"01",
"10",
"10",
"11",
"01",
"01",
"10",
"01",
"10",
"00",
"00",
"01",
"01",
"00",
"11",
"01",
"10",
"10",
"01",
"10",
"11",
"00",
"11",
"00",
"11",
"10",
"01",
"00",
"10",
"00",
"10",
"00",
"00",
"11",
"10",
"01",
"10",
"10",
"10",
"01",
"11",
"10",
"11",
"11",
"11",
"00",
"01",
"01",
"01",
"01",
"01",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"11",
"01",
"11",
"01",
"11",
"11",
"11",
"11",
"11",
"00",
"10",
"10",
"01",
"00",
"11",
"11",
"11",
"11",
"10",
"00",
"00",
"00",
"01",
"00",
"01",
"11",
"11",
"00",
"11",
"11",
"01",
"01",
"11",
"11",
"01",
"01",
"11",
"11",
"11",
"01",
"11",
"10",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"00",
"10",
"10",
"10",
"01",
"01",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"11",
"10",
"10",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"01",
"10",
"00",
"11",
"10",
"10",
"11",
"10",
"10",
"10",
"11",
"00",
"10",
"11",
"00",
"01",
"01",
"00",
"11",
"00",
"00",
"10",
"11",
"11",
"11",
"11",
"00",
"10",
"00",
"00",
"01",
"01",
"01",
"00",
"00",
"01",
"10",
"00",
"10",
"00",
"10",
"01",
"10",
"10",
"00",
"01",
"00",
"11",
"11",
"10",
"11",
"00",
"01",
"11",
"00",
"00",
"01",
"11",
"10",
"10",
"01",
"00",
"01",
"11",
"01",
"01",
"11",
"00",
"00",
"01",
"01",
"00",
"01",
"00",
"01",
"10",
"10",
"00",
"00",
"00",
"11",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",
"00",

others => (others => '0')

);    
begin

process(clk)  begin
	if rising_edge(clk)  then
		if Rd = '1' then
			Data <= rom(conv_integer(addr));  -- First register
		end if;
	end if;
end process;
end Behavioral;


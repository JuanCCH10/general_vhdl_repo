----------------------------------------------------------------------------------
-- Company: SEMAR
-- Engineer: TTE.FRAG.SIA.ELCO. GUILLERMO VICENCIO GUTIERREZ
-- 
-- Create Date:    12:27:30 01/03/2012 
-- Design Name:   MEMORIA
-- Module Name:    RAM_PRF - Behavioral 
-- Project Name: 
-- Target Devices: XC4VSX35-10FF668
-- Tool versions: ISE 13.1
-- Description: ALMACENAR EN EL FPGA LOS DATOS CORRESPONDIENTES A LOS NIVELES
-- DE UNA SE�AL DE FERFIL DE RANGO, ESTA SE�AL FUE MUESTREADA CON EL OSCILOSCOPIO
-- DE UN RADAR BME
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ROM_Mult_alfa is
    generic(Addrbits		: integer;
			DataBits		: integer
				);
	 Port (	Clk : in  STD_LOGIC;
			Addr: in  STD_LOGIC_VECTOR (Addrbits-1 downto 0);
			Rd	: in  STD_LOGIC;
			Data: out  STD_LOGIC_VECTOR (DataBits-1 downto 0));
end ROM_Mult_alfa;

architecture Behavioral of ROM_Mult_alfa is

--ROM PARA GUARDAR LOS comandos para el display oled
TYPE ROM_TYPE IS ARRAY (0 TO 2**Addrbits - 1) OF STD_LOGIC_VECTOR(DATA'range);
SIGNAL ROM: ROM_TYPE := (
--33=>"00001",
--34=>"00010",
--36=>"00100",
--40=>"01000",
--48=>"10000",
--37=>"00101",
--42=>"01010",
--52=>"10100",
--45=>"01101",
--58=>"11010",
--49=>"10001",
--39=>"00111",
--46=>"01110",
--60=>"11100",
--61=>"11101",
--63=>"11111",
--59=>"11011",
--51=>"10011",
--35=>"00011",
--38=>"00110",
--44=>"01100",
--56=>"11000",
--53=>"10101",
--47=>"01111",
--62=>"11110",
--57=>"11001",
--55=>"10111",
--43=>"01011",
--54=>"10110",
--41=>"01001",
--50=>"10010",
----33=>"00001",
--65=>"00010",
--66=>"00100",
--68=>"01000",
--72=>"10000",
--80=>"00101",
--69=>"01010",
--74=>"10100",
--84=>"01101",
--77=>"11010",
--90=>"10001",
--81=>"00111",
--71=>"01110",
--78=>"11100",
--92=>"11101",
--93=>"11111",
--95=>"11011",
--91=>"10011",
--83=>"00011",
--67=>"00110",
--70=>"01100",
--76=>"11000",
--88=>"10101",
--85=>"01111",
--79=>"11110",
--94=>"11001",
--89=>"10111",
--87=>"01011",
--75=>"10110",
--86=>"01001",
--73=>"10010",
--82=>"00001",
----65=>"00010",
--129=>"00100",
--130=>"01000",
--132=>"10000",
--136=>"00101",
--144=>"01010",
--133=>"10100",
--138=>"01101",
--148=>"11010",
--141=>"10001",
--154=>"00111",
--145=>"01110",
--135=>"11100",
--142=>"11101",
--156=>"11111",
--157=>"11011",
--159=>"10011",
--155=>"00011",
--147=>"00110",
--131=>"01100",
--134=>"11000",
--140=>"10101",
--152=>"01111",
--149=>"11110",
--143=>"11001",
--158=>"10111",
--153=>"01011",
--151=>"10110",
--139=>"01001",
--150=>"10010",
--137=>"00001",
--146=>"00010",
----129=>"00100",
--257=>"01000",
--258=>"10000",
--260=>"00101",
--264=>"01010",
--272=>"10100",
--261=>"01101",
--266=>"11010",
--276=>"10001",
--269=>"00111",
--282=>"01110",
--273=>"11100",
--263=>"11101",
--270=>"11111",
--284=>"11011",
--285=>"10011",
--287=>"00011",
--283=>"00110",
--275=>"01100",
--259=>"11000",
--262=>"10101",
--268=>"01111",
--280=>"11110",
--277=>"11001",
--271=>"10111",
--286=>"01011",
--281=>"10110",
--279=>"01001",
--267=>"10010",
--278=>"00001",
--265=>"00010",
--274=>"00100",
----257=>"01000",
--513=>"10000",
--514=>"00101",
--516=>"01010",
--520=>"10100",
--528=>"01101",
--517=>"11010",
--522=>"10001",
--532=>"00111",
--525=>"01110",
--538=>"11100",
--529=>"11101",
--519=>"11111",
--526=>"11011",
--540=>"10011",
--541=>"00011",
--543=>"00110",
--539=>"01100",
--531=>"11000",
--515=>"10101",
--518=>"01111",
--524=>"11110",
--536=>"11001",
--533=>"10111",
--527=>"01011",
--542=>"10110",
--537=>"01001",
--535=>"10010",
--523=>"00001",
--534=>"00010",
--521=>"00100",
--530=>"01000",
----513=>"10000",
--161=>"00101",
--162=>"01010",
--164=>"10100",
--168=>"01101",
--176=>"11010",
--165=>"10001",
--170=>"00111",
--180=>"01110",
--173=>"11100",
--186=>"11101",
--177=>"11111",
--167=>"11011",
--174=>"10011",
--188=>"00011",
--189=>"00110",
--191=>"01100",
--187=>"11000",
--179=>"10101",
--163=>"01111",
--166=>"11110",
--172=>"11001",
--184=>"10111",
--181=>"01011",
--175=>"10110",
--190=>"01001",
--185=>"10010",
--183=>"00001",
--171=>"00010",
--182=>"00100",
--169=>"01000",
--178=>"10000",
----161=>"00101",
--321=>"01010",
--322=>"10100",
--324=>"01101",
--328=>"11010",
--336=>"10001",
--325=>"00111",
--330=>"01110",
--340=>"11100",
--333=>"11101",
--346=>"11111",
--337=>"11011",
--327=>"10011",
--334=>"00011",
--348=>"00110",
--349=>"01100",
--351=>"11000",
--347=>"10101",
--339=>"01111",
--323=>"11110",
--326=>"11001",
--332=>"10111",
--344=>"01011",
--341=>"10110",
--335=>"01001",
--350=>"10010",
--345=>"00001",
--343=>"00010",
--331=>"00100",
--342=>"01000",
--329=>"10000",
--338=>"00101",
----321=>"01010",
--641=>"10100",
--642=>"01101",
--644=>"11010",
--648=>"10001",
--656=>"00111",
--645=>"01110",
--650=>"11100",
--660=>"11101",
--653=>"11111",
--666=>"11011",
--657=>"10011",
--647=>"00011",
--654=>"00110",
--668=>"01100",
--669=>"11000",
--671=>"10101",
--667=>"01111",
--659=>"11110",
--643=>"11001",
--646=>"10111",
--652=>"01011",
--664=>"10110",
--661=>"01001",
--655=>"10010",
--670=>"00001",
--665=>"00010",
--663=>"00100",
--651=>"01000",
--662=>"10000",
--649=>"00101",
--658=>"01010",
----641=>"10100",
--417=>"01101",
--418=>"11010",
--420=>"10001",
--424=>"00111",
--432=>"01110",
--421=>"11100",
--426=>"11101",
--436=>"11111",
--429=>"11011",
--442=>"10011",
--433=>"00011",
--423=>"00110",
--430=>"01100",
--444=>"11000",
--445=>"10101",
--447=>"01111",
--443=>"11110",
--435=>"11001",
--419=>"10111",
--422=>"01011",
--428=>"10110",
--440=>"01001",
--437=>"10010",
--431=>"00001",
--446=>"00010",
--441=>"00100",
--439=>"01000",
--427=>"10000",
--438=>"00101",
--425=>"01010",
--434=>"10100",
----417=>"01101",
--833=>"11010",
--834=>"10001",
--836=>"00111",
--840=>"01110",
--848=>"11100",
--837=>"11101",
--842=>"11111",
--852=>"11011",
--845=>"10011",
--858=>"00011",
--849=>"00110",
--839=>"01100",
--846=>"11000",
--860=>"10101",
--861=>"01111",
--863=>"11110",
--859=>"11001",
--851=>"10111",
--835=>"01011",
--838=>"10110",
--844=>"01001",
--856=>"10010",
--853=>"00001",
--847=>"00010",
--862=>"00100",
--857=>"01000",
--855=>"10000",
--843=>"00101",
--854=>"01010",
--841=>"10100",
--850=>"01101",
----833=>"11010",
--545=>"10001",
--546=>"00111",
--548=>"01110",
--552=>"11100",
--560=>"11101",
--549=>"11111",
--554=>"11011",
--564=>"10011",
--557=>"00011",
--570=>"00110",
--561=>"01100",
--551=>"11000",
--558=>"10101",
--572=>"01111",
--573=>"11110",
--575=>"11001",
--571=>"10111",
--563=>"01011",
--547=>"10110",
--550=>"01001",
--556=>"10010",
--568=>"00001",
--565=>"00010",
--559=>"00100",
--574=>"01000",
--569=>"10000",
--567=>"00101",
--555=>"01010",
--566=>"10100",
--553=>"01101",
--562=>"11010",
----545=>"10001",
--225=>"00111",
--226=>"01110",
--228=>"11100",
--232=>"11101",
--240=>"11111",
--229=>"11011",
--234=>"10011",
--244=>"00011",
--237=>"00110",
--250=>"01100",
--241=>"11000",
--231=>"10101",
--238=>"01111",
--252=>"11110",
--253=>"11001",
--255=>"10111",
--251=>"01011",
--243=>"10110",
--227=>"01001",
--230=>"10010",
--236=>"00001",
--248=>"00010",
--245=>"00100",
--239=>"01000",
--254=>"10000",
--249=>"00101",
--247=>"01010",
--235=>"10100",
--246=>"01101",
--233=>"11010",
--242=>"10001",
----225=>"00111",
--449=>"01110",
--450=>"11100",
--452=>"11101",
--456=>"11111",
--464=>"11011",
--453=>"10011",
--458=>"00011",
--468=>"00110",
--461=>"01100",
--474=>"11000",
--465=>"10101",
--455=>"01111",
--462=>"11110",
--476=>"11001",
--477=>"10111",
--479=>"01011",
--475=>"10110",
--467=>"01001",
--451=>"10010",
--454=>"00001",
--460=>"00010",
--472=>"00100",
--469=>"01000",
--463=>"10000",
--478=>"00101",
--473=>"01010",
--471=>"10100",
--459=>"01101",
--470=>"11010",
--457=>"10001",
--466=>"00111",
----449=>"01110",
--897=>"11100",
--898=>"11101",
--900=>"11111",
--904=>"11011",
--912=>"10011",
--901=>"00011",
--906=>"00110",
--916=>"01100",
--909=>"11000",
--922=>"10101",
--913=>"01111",
--903=>"11110",
--910=>"11001",
--924=>"10111",
--925=>"01011",
--927=>"10110",
--923=>"01001",
--915=>"10010",
--899=>"00001",
--902=>"00010",
--908=>"00100",
--920=>"01000",
--917=>"10000",
--911=>"00101",
--926=>"01010",
--921=>"10100",
--919=>"01101",
--907=>"11010",
--918=>"10001",
--905=>"00111",
--914=>"01110",
----897=>"11100",
--929=>"11101",
--930=>"11111",
--932=>"11011",
--936=>"10011",
--944=>"00011",
--933=>"00110",
--938=>"01100",
--948=>"11000",
--941=>"10101",
--954=>"01111",
--945=>"11110",
--935=>"11001",
--942=>"10111",
--956=>"01011",
--957=>"10110",
--959=>"01001",
--955=>"10010",
--947=>"00001",
--931=>"00010",
--934=>"00100",
--940=>"01000",
--952=>"10000",
--949=>"00101",
--943=>"01010",
--958=>"10100",
--953=>"01101",
--951=>"11010",
--939=>"10001",
--950=>"00111",
--937=>"01110",
--946=>"11100",
----929=>"11101",
--993=>"11111",
--994=>"11011",
--996=>"10011",
--1000=>"00011",
--1008=>"00110",
--997=>"01100",
--1002=>"11000",
--1012=>"10101",
--1005=>"01111",
--1018=>"11110",
--1009=>"11001",
--999=>"10111",
--1006=>"01011",
--1020=>"10110",
--1021=>"01001",
--1023=>"10010",
--1019=>"00001",
--1011=>"00010",
--995=>"00100",
--998=>"01000",
--1004=>"10000",
--1016=>"00101",
--1013=>"01010",
--1007=>"10100",
--1022=>"01101",
--1017=>"11010",
--1015=>"10001",
--1003=>"00111",
--1014=>"01110",
--1001=>"11100",
--1010=>"11101",
----993=>"11111",
--865=>"11011",
--866=>"10011",
--868=>"00011",
--872=>"00110",
--880=>"01100",
--869=>"11000",
--874=>"10101",
--884=>"01111",
--877=>"11110",
--890=>"11001",
--881=>"10111",
--871=>"01011",
--878=>"10110",
--892=>"01001",
--893=>"10010",
--895=>"00001",
--891=>"00010",
--883=>"00100",
--867=>"01000",
--870=>"10000",
--876=>"00101",
--888=>"01010",
--885=>"10100",
--879=>"01101",
--894=>"11010",
--889=>"10001",
--887=>"00111",
--875=>"01110",
--886=>"11100",
--873=>"11101",
--882=>"11111",
----865=>"11011",
--609=>"10011",
--610=>"00011",
--612=>"00110",
--616=>"01100",
--624=>"11000",
--613=>"10101",
--618=>"01111",
--628=>"11110",
--621=>"11001",
--634=>"10111",
--625=>"01011",
--615=>"10110",
--622=>"01001",
--636=>"10010",
--637=>"00001",
--639=>"00010",
--635=>"00100",
--627=>"01000",
--611=>"10000",
--614=>"00101",
--620=>"01010",
--632=>"10100",
--629=>"01101",
--623=>"11010",
--638=>"10001",
--633=>"00111",
--631=>"01110",
--619=>"11100",
--630=>"11101",
--617=>"11111",
--626=>"11011",
----609=>"10011",
--97=>"00011",
--98=>"00110",
--100=>"01100",
--104=>"11000",
--112=>"10101",
--101=>"01111",
--106=>"11110",
--116=>"11001",
--109=>"10111",
--122=>"01011",
--113=>"10110",
--103=>"01001",
--110=>"10010",
--124=>"00001",
--125=>"00010",
--127=>"00100",
--123=>"01000",
--115=>"10000",
--99=>"00101",
--102=>"01010",
--108=>"10100",
--120=>"01101",
--117=>"11010",
--111=>"10001",
--126=>"00111",
--121=>"01110",
--119=>"11100",
--107=>"11101",
--118=>"11111",
--105=>"11011",
--114=>"10011",
----97=>"00011",
--193=>"00110",
--194=>"01100",
--196=>"11000",
--200=>"10101",
--208=>"01111",
--197=>"11110",
--202=>"11001",
--212=>"10111",
--205=>"01011",
--218=>"10110",
--209=>"01001",
--199=>"10010",
--206=>"00001",
--220=>"00010",
--221=>"00100",
--223=>"01000",
--219=>"10000",
--211=>"00101",
--195=>"01010",
--198=>"10100",
--204=>"01101",
--216=>"11010",
--213=>"10001",
--207=>"00111",
--222=>"01110",
--217=>"11100",
--215=>"11101",
--203=>"11111",
--214=>"11011",
--201=>"10011",
--210=>"00011",
----193=>"00110",
--385=>"01100",
--386=>"11000",
--388=>"10101",
--392=>"01111",
--400=>"11110",
--389=>"11001",
--394=>"10111",
--404=>"01011",
--397=>"10110",
--410=>"01001",
--401=>"10010",
--391=>"00001",
--398=>"00010",
--412=>"00100",
--413=>"01000",
--415=>"10000",
--411=>"00101",
--403=>"01010",
--387=>"10100",
--390=>"01101",
--396=>"11010",
--408=>"10001",
--405=>"00111",
--399=>"01110",
--414=>"11100",
--409=>"11101",
--407=>"11111",
--395=>"11011",
--406=>"10011",
--393=>"00011",
--402=>"00110",
----385=>"01100",
--769=>"11000",
--770=>"10101",
--772=>"01111",
--776=>"11110",
--784=>"11001",
--773=>"10111",
--778=>"01011",
--788=>"10110",
--781=>"01001",
--794=>"10010",
--785=>"00001",
--775=>"00010",
--782=>"00100",
--796=>"01000",
--797=>"10000",
--799=>"00101",
--795=>"01010",
--787=>"10100",
--771=>"01101",
--774=>"11010",
--780=>"10001",
--792=>"00111",
--789=>"01110",
--783=>"11100",
--798=>"11101",
--793=>"11111",
--791=>"11011",
--779=>"10011",
--790=>"00011",
--777=>"00110",
--786=>"01100",
----769=>"11000",
--673=>"10101",
--674=>"01111",
--676=>"11110",
--680=>"11001",
--688=>"10111",
--677=>"01011",
--682=>"10110",
--692=>"01001",
--685=>"10010",
--698=>"00001",
--689=>"00010",
--679=>"00100",
--686=>"01000",
--700=>"10000",
--701=>"00101",
--703=>"01010",
--699=>"10100",
--691=>"01101",
--675=>"11010",
--678=>"10001",
--684=>"00111",
--696=>"01110",
--693=>"11100",
--687=>"11101",
--702=>"11111",
--697=>"11011",
--695=>"10011",
--683=>"00011",
--694=>"00110",
--681=>"01100",
--690=>"11000",
----673=>"10101",
--481=>"01111",
--482=>"11110",
--484=>"11001",
--488=>"10111",
--496=>"01011",
--485=>"10110",
--490=>"01001",
--500=>"10010",
--493=>"00001",
--506=>"00010",
--497=>"00100",
--487=>"01000",
--494=>"10000",
--508=>"00101",
--509=>"01010",
--511=>"10100",
--507=>"01101",
--499=>"11010",
--483=>"10001",
--486=>"00111",
--492=>"01110",
--504=>"11100",
--501=>"11101",
--495=>"11111",
--510=>"11011",
--505=>"10011",
--503=>"00011",
--491=>"00110",
--502=>"01100",
--489=>"11000",
--498=>"10101",
----481=>"01111",
--961=>"11110",
--962=>"11001",
--964=>"10111",
--968=>"01011",
--976=>"10110",
--965=>"01001",
--970=>"10010",
--980=>"00001",
--973=>"00010",
--986=>"00100",
--977=>"01000",
--967=>"10000",
--974=>"00101",
--988=>"01010",
--989=>"10100",
--991=>"01101",
--987=>"11010",
--979=>"10001",
--963=>"00111",
--966=>"01110",
--972=>"11100",
--984=>"11101",
--981=>"11111",
--975=>"11011",
--990=>"10011",
--985=>"00011",
--983=>"00110",
--971=>"01100",
--982=>"11000",
--969=>"10101",
--978=>"01111",
----961=>"11110",
--801=>"11001",
--802=>"10111",
--804=>"01011",
--808=>"10110",
--816=>"01001",
--805=>"10010",
--810=>"00001",
--820=>"00010",
--813=>"00100",
--826=>"01000",
--817=>"10000",
--807=>"00101",
--814=>"01010",
--828=>"10100",
--829=>"01101",
--831=>"11010",
--827=>"10001",
--819=>"00111",
--803=>"01110",
--806=>"11100",
--812=>"11101",
--824=>"11111",
--821=>"11011",
--815=>"10011",
--830=>"00011",
--825=>"00110",
--823=>"01100",
--811=>"11000",
--822=>"10101",
--809=>"01111",
--818=>"11110",
----801=>"11001",
--737=>"10111",
--738=>"01011",
--740=>"10110",
--744=>"01001",
--752=>"10010",
--741=>"00001",
--746=>"00010",
--756=>"00100",
--749=>"01000",
--762=>"10000",
--753=>"00101",
--743=>"01010",
--750=>"10100",
--764=>"01101",
--765=>"11010",
--767=>"10001",
--763=>"00111",
--755=>"01110",
--739=>"11100",
--742=>"11101",
--748=>"11111",
--760=>"11011",
--757=>"10011",
--751=>"00011",
--766=>"00110",
--761=>"01100",
--759=>"11000",
--747=>"10101",
--758=>"01111",
--745=>"11110",
--754=>"11001",
----737=>"10111",
--353=>"01011",
--354=>"10110",
--356=>"01001",
--360=>"10010",
--368=>"00001",
--357=>"00010",
--362=>"00100",
--372=>"01000",
--365=>"10000",
--378=>"00101",
--369=>"01010",
--359=>"10100",
--366=>"01101",
--380=>"11010",
--381=>"10001",
--383=>"00111",
--379=>"01110",
--371=>"11100",
--355=>"11101",
--358=>"11111",
--364=>"11011",
--376=>"10011",
--373=>"00011",
--367=>"00110",
--382=>"01100",
--377=>"11000",
--375=>"10101",
--363=>"01111",
--374=>"11110",
--361=>"11001",
--370=>"10111",
----353=>"01011",
--705=>"10110",
--706=>"01001",
--708=>"10010",
--712=>"00001",
--720=>"00010",
--709=>"00100",
--714=>"01000",
--724=>"10000",
--717=>"00101",
--730=>"01010",
--721=>"10100",
--711=>"01101",
--718=>"11010",
--732=>"10001",
--733=>"00111",
--735=>"01110",
--731=>"11100",
--723=>"11101",
--707=>"11111",
--710=>"11011",
--716=>"10011",
--728=>"00011",
--725=>"00110",
--719=>"01100",
--734=>"11000",
--729=>"10101",
--727=>"01111",
--715=>"11110",
--726=>"11001",
--713=>"10111",
--722=>"01011",
----705=>"10110",
--289=>"01001",
--290=>"10010",
--292=>"00001",
--296=>"00010",
--304=>"00100",
--293=>"01000",
--298=>"10000",
--308=>"00101",
--301=>"01010",
--314=>"10100",
--305=>"01101",
--295=>"11010",
--302=>"10001",
--316=>"00111",
--317=>"01110",
--319=>"11100",
--315=>"11101",
--307=>"11111",
--291=>"11011",
--294=>"10011",
--300=>"00011",
--312=>"00110",
--309=>"01100",
--303=>"11000",
--318=>"10101",
--313=>"01111",
--311=>"11110",
--299=>"11001",
--310=>"10111",
--297=>"01011",
--306=>"10110",
----289=>"01001",
--577=>"10010",
--578=>"00001",
--580=>"00010",
--584=>"00100",
--592=>"01000",
--581=>"10000",
--586=>"00101",
--596=>"01010",
--589=>"10100",
--602=>"01101",
--593=>"11010",
--583=>"10001",
--590=>"00111",
--604=>"01110",
--605=>"11100",
--607=>"11101",
--603=>"11111",
--595=>"11011",
--579=>"10011",
--582=>"00011",
--588=>"00110",
--600=>"01100",
--597=>"11000",
--591=>"10101",
--606=>"01111",
--601=>"11110",
--599=>"11001",
--587=>"10111",
--598=>"01011",
--585=>"10110",
--594=>"01001",


----577=>"10010",
----33=>"00001",
----34=>"00010",
----36=>"00100",
----40=>"01000",
----48=>"10000",
----37=>"00101",
----42=>"01010",
----52=>"10100",
----45=>"01101",
----58=>"11010",
----49=>"10001",
----39=>"00111",
----46=>"01110",
----60=>"11100",
----61=>"11101",
----63=>"11111",
----59=>"11011",
----51=>"10011",
----35=>"00011",
----38=>"00110",
----44=>"01100",
----56=>"11000",
----53=>"10101",
----47=>"01111",
----62=>"11110",
----57=>"11001",
----55=>"10111",
----43=>"01011",
----54=>"10110",
----41=>"01001",
----50=>"10010",
----33=>"00001",

65 => "000001",
66 => "000010",
68 => "000100",
72 => "001000",
80 => "010000",
96 => "100000",
67 => "000011",
70 => "000110",
76 => "001100",
88 => "011000",
112=> "110000",
99 => "100011",
69 => "000101",
74 => "001010",
84 => "010100",
104=> "101000",
83 => "010011",
102=> "100110",
79 => "001111",
94 => "011110",
124=> "111100",
123=> "111011",
117=> "110101",
105=> "101001",
81 => "010001",
98 => "100010",
71 => "000111",
78 => "001110",
92 => "011100",
120=> "111000",
115=> "110011",
101=> "100101",
73 => "001001",
82 => "010010",
100=> "100100",
75 => "001011",
86 => "010110",
108=> "101100",
91 => "011011",
118=> "110110",
111=> "101111",
93 => "011101",
122=> "111010",
119=> "110111",
109=> "101101",
89 => "011001",
114=> "110010",
103=> "100111",
77 => "001101",
90 => "011010",
116=> "110100",
107=> "101011",
85 => "010101",
106=> "101010",
87 => "010111",
110=> "101110",
95 => "011111",
126=> "111110",
127=> "111111",
125=> "111101",
121=> "111001",
113=> "110001",
97 => "100001",
   
129=> "000010",
130=> "000100",
132=> "001000",
136=> "010000",
144=> "100000",
160=> "000011",
131=> "000110",
134=> "001100",
140=> "011000",
152=> "110000",
176=> "100011",
163=> "000101",
133=> "001010",
138=> "010100",
148=> "101000",
168=> "010011",
147=> "100110",
166=> "001111",
143=> "011110",
158=> "111100",
188=> "111011",
187=> "110101",
181=> "101001",
169=> "010001",
145=> "100010",
162=> "000111",
135=> "001110",
142=> "011100",
156=> "111000",
184=> "110011",
179=> "100101",
165=> "001001",
137=> "010010",
146=> "100100",
164=> "001011",
139=> "010110",
150=> "101100",
172=> "011011",
155=> "110110",
182=> "101111",
175=> "011101",
157=> "111010",
186=> "110111",
183=> "101101",
173=> "011001",
153=> "110010",
178=> "100111",
167=> "001101",
141=> "011010",
154=> "110100",
180=> "101011",
171=> "010101",
149=> "101010",
170=> "010111",
151=> "101110",
174=> "011111",
159=> "111110",
190=> "111111",
191=> "111101",
189=> "111001",
185=> "110001",
177=> "100001",
161=> "000001",

257=> "000100",
258=> "001000",
260=> "010000",
264=> "100000",
272=> "000011",
288=> "000110",
259=> "001100",
262=> "011000",
268=> "110000",
280=> "100011",
304=> "000101",
291=> "001010",
261=> "010100",
266=> "101000",
276=> "010011",
296=> "100110",
275=> "001111",
294=> "011110",
271=> "111100",
286=> "111011",
316=> "110101",
315=> "101001",
309=> "010001",
297=> "100010",
273=> "000111",
290=> "001110",
263=> "011100",
270=> "111000",
284=> "110011",
312=> "100101",
307=> "001001",
293=> "010010",
265=> "100100",
274=> "001011",
292=> "010110",
267=> "101100",
278=> "011011",
300=> "110110",
283=> "101111",
310=> "011101",
303=> "111010",
285=> "110111",
314=> "101101",
311=> "011001",
301=> "110010",
281=> "100111",
306=> "001101",
295=> "011010",
269=> "110100",
282=> "101011",
308=> "010101",
299=> "101010",
277=> "010111",
298=> "101110",
279=> "011111",
302=> "111110",
287=> "111111",
318=> "111101",
319=> "111001",
317=> "110001",
313=> "100001",
305=> "000001",
289=> "000010",

513=> "001000",
514=> "010000",
516=> "100000",
520=> "000011",
528=> "000110",
544=> "001100",
515=> "011000",
518=> "110000",
524=> "100011",
536=> "000101",
560=> "001010",
547=> "010100",
517=> "101000",
522=> "010011",
532=> "100110",
552=> "001111",
531=> "011110",
550=> "111100",
527=> "111011",
542=> "110101",
572=> "101001",
571=> "010001",
565=> "100010",
553=> "000111",
529=> "001110",
546=> "011100",
519=> "111000",
526=> "110011",
540=> "100101",
568=> "001001",
563=> "010010",
549=> "100100",
521=> "001011",
530=> "010110",
548=> "101100",
523=> "011011",
534=> "110110",
556=> "101111",
539=> "011101",
566=> "111010",
559=> "110111",
541=> "101101",
570=> "011001",
567=> "110010",
557=> "100111",
537=> "001101",
562=> "011010",
551=> "110100",
525=> "101011",
538=> "010101",
564=> "101010",
555=> "010111",
533=> "101110",
554=> "011111",
535=> "111110",
558=> "111111",
543=> "111101",
574=> "111001",
575=> "110001",
573=> "100001",
569=> "000001",
561=> "000010",
545=> "000100",

1025=>"010000",
1026=>"100000",
1028=>"000011",
1032=>"000110",
1040=>"001100",
1056=>"011000",
1027=>"110000",
1030=>"100011",
1036=>"000101",
1048=>"001010",
1072=>"010100",
1059=>"101000",
1029=>"010011",
1034=>"100110",
1044=>"001111",
1064=>"011110",
1043=>"111100",
1062=>"111011",
1039=>"110101",
1054=>"101001",
1084=>"010001",
1083=>"100010",
1077=>"000111",
1065=>"001110",
1041=>"011100",
1058=>"111000",
1031=>"110011",
1038=>"100101",
1052=>"001001",
1080=>"010010",
1075=>"100100",
1061=>"001011",
1033=>"010110",
1042=>"101100",
1060=>"011011",
1035=>"110110",
1046=>"101111",
1068=>"011101",
1051=>"111010",
1078=>"110111",
1071=>"101101",
1053=>"011001",
1082=>"110010",
1079=>"100111",
1069=>"001101",
1049=>"011010",
1074=>"110100",
1063=>"101011",
1037=>"010101",
1050=>"101010",
1076=>"010111",
1067=>"101110",
1045=>"011111",
1066=>"111110",
1047=>"111111",
1070=>"111101",
1055=>"111001",
1086=>"110001",
1087=>"100001",
1085=>"000001",
1081=>"000010",
1073=>"000100",
1057=>"001000",

2049=>"100000",
2050=>"000011",
2052=>"000110",
2056=>"001100",
2064=>"011000",
2080=>"110000",
2051=>"100011",
2054=>"000101",
2060=>"001010",
2072=>"010100",
2096=>"101000",
2083=>"010011",
2053=>"100110",
2058=>"001111",
2068=>"011110",
2088=>"111100",
2067=>"111011",
2086=>"110101",
2063=>"101001",
2078=>"010001",
2108=>"100010",
2107=>"000111",
2101=>"001110",
2089=>"011100",
2065=>"111000",
2082=>"110011",
2055=>"100101",
2062=>"001001",
2076=>"010010",
2104=>"100100",
2099=>"001011",
2085=>"010110",
2057=>"101100",
2066=>"011011",
2084=>"110110",
2059=>"101111",
2070=>"011101",
2092=>"111010",
2075=>"110111",
2102=>"101101",
2095=>"011001",
2077=>"110010",
2106=>"100111",
2103=>"001101",
2093=>"011010",
2073=>"110100",
2098=>"101011",
2087=>"010101",
2061=>"101010",
2074=>"010111",
2100=>"101110",
2091=>"011111",
2069=>"111110",
2090=>"111111",
2071=>"111101",
2094=>"111001",
2079=>"110001",
2110=>"100001",
2111=>"000001",
2109=>"000010",
2105=>"000100",
2097=>"001000",
2081=>"010000",

193 =>"000011",
194 =>"000110",
196 =>"001100",
200 =>"011000",
208 =>"110000",
224 =>"100011",
195 =>"000101",
198 =>"001010",
204 =>"010100",
216 =>"101000",
240 =>"010011",
227 =>"100110",
197 =>"001111",
202 =>"011110",
212 =>"111100",
232 =>"111011",
211 =>"110101",
230 =>"101001",
207 =>"010001",
222 =>"100010",
252 =>"000111",
251 =>"001110",
245 =>"011100",
233 =>"111000",
209 =>"110011",
226 =>"100101",
199 =>"001001",
206 =>"010010",
220 =>"100100",
248 =>"001011",
243 =>"010110",
229 =>"101100",
201 =>"011011",
210 =>"110110",
228 =>"101111",
203 =>"011101",
214 =>"111010",
236 =>"110111",
219 =>"101101",
246 =>"011001",
239 =>"110010",
221 =>"100111",
250 =>"001101",
247 =>"011010",
237 =>"110100",
217 =>"101011",
242 =>"010101",
231 =>"101010",
205 =>"010111",
218 =>"101110",
244 =>"011111",
235 =>"111110",
213 =>"111111",
234 =>"111101",
215 =>"111001",
238 =>"110001",
223 =>"100001",
254 =>"000001",
255 =>"000010",
253 =>"000100",
249 =>"001000",
241 =>"010000",
225 =>"100000",

385 =>"000110",
386 =>"001100",
388 =>"011000",
392 =>"110000",
400 =>"100011",
416 =>"000101",
387 =>"001010",
390 =>"010100",
396 =>"101000",
408 =>"010011",
432 =>"100110",
419 =>"001111",
389 =>"011110",
394 =>"111100",
404 =>"111011",
424 =>"110101",
403 =>"101001",
422 =>"010001",
399 =>"100010",
414 =>"000111",
444 =>"001110",
443 =>"011100",
437 =>"111000",
425 =>"110011",
401 =>"100101",
418 =>"001001",
391 =>"010010",
398 =>"100100",
412 =>"001011",
440 =>"010110",
435 =>"101100",
421 =>"011011",
393 =>"110110",
402 =>"101111",
420 =>"011101",
395 =>"111010",
406 =>"110111",
428 =>"101101",
411 =>"011001",
438 =>"110010",
431 =>"100111",
413 =>"001101",
442 =>"011010",
439 =>"110100",
429 =>"101011",
409 =>"010101",
434 =>"101010",
423 =>"010111",
397 =>"101110",
410 =>"011111",
436 =>"111110",
427 =>"111111",
405 =>"111101",
426 =>"111001",
407 =>"110001",
430 =>"100001",
415 =>"000001",
446 =>"000010",
447 =>"000100",
445 =>"001000",
441 =>"010000",
433 =>"100000",
417 =>"000011",
      
769 =>"001100",
770 =>"011000",
772 =>"110000",
776 =>"100011",
784 =>"000101",
800 =>"001010",
771 =>"010100",
774 =>"101000",
780 =>"010011",
792 =>"100110",
816 =>"001111",
803 =>"011110",
773 =>"111100",
778 =>"111011",
788 =>"110101",
808 =>"101001",
787 =>"010001",
806 =>"100010",
783 =>"000111",
798 =>"001110",
828 =>"011100",
827 =>"111000",
821 =>"110011",
809 =>"100101",
785 =>"001001",
802 =>"010010",
775 =>"100100",
782 =>"001011",
796 =>"010110",
824 =>"101100",
819 =>"011011",
805 =>"110110",
777 =>"101111",
786 =>"011101",
804 =>"111010",
779 =>"110111",
790 =>"101101",
812 =>"011001",
795 =>"110010",
822 =>"100111",
815 =>"001101",
797 =>"011010",
826 =>"110100",
823 =>"101011",
813 =>"010101",
793 =>"101010",
818 =>"010111",
807 =>"101110",
781 =>"011111",
794 =>"111110",
820 =>"111111",
811 =>"111101",
789 =>"111001",
810 =>"110001",
791 =>"100001",
814 =>"000001",
799 =>"000010",
830 =>"000100",
831 =>"001000",
829 =>"010000",
825 =>"100000",
817 =>"000011",
801 =>"000110",
      
1537=>"011000",
1538=>"110000",
1540=>"100011",
1544=>"000101",
1552=>"001010",
1568=>"010100",
1539=>"101000",
1542=>"010011",
1548=>"100110",
1560=>"001111",
1584=>"011110",
1571=>"111100",
1541=>"111011",
1546=>"110101",
1556=>"101001",
1576=>"010001",
1555=>"100010",
1574=>"000111",
1551=>"001110",
1566=>"011100",
1596=>"111000",
1595=>"110011",
1589=>"100101",
1577=>"001001",
1553=>"010010",
1570=>"100100",
1543=>"001011",
1550=>"010110",
1564=>"101100",
1592=>"011011",
1587=>"110110",
1573=>"101111",
1545=>"011101",
1554=>"111010",
1572=>"110111",
1547=>"101101",
1558=>"011001",
1580=>"110010",
1563=>"100111",
1590=>"001101",
1583=>"011010",
1565=>"110100",
1594=>"101011",
1591=>"010101",
1581=>"101010",
1561=>"010111",
1586=>"101110",
1575=>"011111",
1549=>"111110",
1562=>"111111",
1588=>"111101",
1579=>"111001",
1557=>"110001",
1578=>"100001",
1559=>"000001",
1582=>"000010",
1567=>"000100",
1598=>"001000",
1599=>"010000",
1597=>"100000",
1593=>"000011",
1585=>"000110",
1569=>"001100",
      
3073=>"110000",
3074=>"100011",
3076=>"000101",
3080=>"001010",
3088=>"010100",
3104=>"101000",
3075=>"010011",
3078=>"100110",
3084=>"001111",
3096=>"011110",
3120=>"111100",
3107=>"111011",
3077=>"110101",
3082=>"101001",
3092=>"010001",
3112=>"100010",
3091=>"000111",
3110=>"001110",
3087=>"011100",
3102=>"111000",
3132=>"110011",
3131=>"100101",
3125=>"001001",
3113=>"010010",
3089=>"100100",
3106=>"001011",
3079=>"010110",
3086=>"101100",
3100=>"011011",
3128=>"110110",
3123=>"101111",
3109=>"011101",
3081=>"111010",
3090=>"110111",
3108=>"101101",
3083=>"011001",
3094=>"110010",
3116=>"100111",
3099=>"001101",
3126=>"011010",
3119=>"110100",
3101=>"101011",
3130=>"010101",
3127=>"101010",
3117=>"010111",
3097=>"101110",
3122=>"011111",
3111=>"111110",
3085=>"111111",
3098=>"111101",
3124=>"111001",
3115=>"110001",
3093=>"100001",
3114=>"000001",
3095=>"000010",
3118=>"000100",
3103=>"001000",
3134=>"010000",
3135=>"100000",
3133=>"000011",
3129=>"000110",
3121=>"001100",
3105=>"011000",
      
2241=>"100011",
2242=>"000101",
2244=>"001010",
2248=>"010100",
2256=>"101000",
2272=>"010011",
2243=>"100110",
2246=>"001111",
2252=>"011110",
2264=>"111100",
2288=>"111011",
2275=>"110101",
2245=>"101001",
2250=>"010001",
2260=>"100010",
2280=>"000111",
2259=>"001110",
2278=>"011100",
2255=>"111000",
2270=>"110011",
2300=>"100101",
2299=>"001001",
2293=>"010010",
2281=>"100100",
2257=>"001011",
2274=>"010110",
2247=>"101100",
2254=>"011011",
2268=>"110110",
2296=>"101111",
2291=>"011101",
2277=>"111010",
2249=>"110111",
2258=>"101101",
2276=>"011001",
2251=>"110010",
2262=>"100111",
2284=>"001101",
2267=>"011010",
2294=>"110100",
2287=>"101011",
2269=>"010101",
2298=>"101010",
2295=>"010111",
2285=>"101110",
2265=>"011111",
2290=>"111110",
2279=>"111111",
2253=>"111101",
2266=>"111001",
2292=>"110001",
2283=>"100001",
2261=>"000001",
2282=>"000010",
2263=>"000100",
2286=>"001000",
2271=>"010000",
2302=>"100000",
2303=>"000011",
2301=>"000110",
2297=>"001100",
2289=>"011000",
2273=>"110000",
      
321 =>"000101",
322 =>"001010",
324 =>"010100",
328 =>"101000",
336 =>"010011",
352 =>"100110",
323 =>"001111",
326 =>"011110",
332 =>"111100",
344 =>"111011",
368 =>"110101",
355 =>"101001",
325 =>"010001",
330 =>"100010",
340 =>"000111",
360 =>"001110",
339 =>"011100",
358 =>"111000",
335 =>"110011",
350 =>"100101",
380 =>"001001",
379 =>"010010",
373 =>"100100",
361 =>"001011",
337 =>"010110",
354 =>"101100",
327 =>"011011",
334 =>"110110",
348 =>"101111",
376 =>"011101",
371 =>"111010",
357 =>"110111",
329 =>"101101",
338 =>"011001",
356 =>"110010",
331 =>"100111",
342 =>"001101",
364 =>"011010",
347 =>"110100",
374 =>"101011",
367 =>"010101",
349 =>"101010",
378 =>"010111",
375 =>"101110",
365 =>"011111",
345 =>"111110",
370 =>"111111",
359 =>"111101",
333 =>"111001",
346 =>"110001",
372 =>"100001",
363 =>"000001",
341 =>"000010",
362 =>"000100",
343 =>"001000",
366 =>"010000",
351 =>"100000",
382 =>"000011",
383 =>"000110",
381 =>"001100",
377 =>"011000",
369 =>"110000",
353 =>"100011",
      
641 =>"001010",
642 =>"010100",
644 =>"101000",
648 =>"010011",
656 =>"100110",
672 =>"001111",
643 =>"011110",
646 =>"111100",
652 =>"111011",
664 =>"110101",
688 =>"101001",
675 =>"010001",
645 =>"100010",
650 =>"000111",
660 =>"001110",
680 =>"011100",
659 =>"111000",
678 =>"110011",
655 =>"100101",
670 =>"001001",
700 =>"010010",
699 =>"100100",
693 =>"001011",
681 =>"010110",
657 =>"101100",
674 =>"011011",
647 =>"110110",
654 =>"101111",
668 =>"011101",
696 =>"111010",
691 =>"110111",
677 =>"101101",
649 =>"011001",
658 =>"110010",
676 =>"100111",
651 =>"001101",
662 =>"011010",
684 =>"110100",
667 =>"101011",
694 =>"010101",
687 =>"101010",
669 =>"010111",
698 =>"101110",
695 =>"011111",
685 =>"111110",
665 =>"111111",
690 =>"111101",
679 =>"111001",
653 =>"110001",
666 =>"100001",
692 =>"000001",
683 =>"000010",
661 =>"000100",
682 =>"001000",
663 =>"010000",
686 =>"100000",
671 =>"000011",
702 =>"000110",
703 =>"001100",
701 =>"011000",
697 =>"110000",
689 =>"100011",
673 =>"000101",
      
1281=>"010100",
1282=>"101000",
1284=>"010011",
1288=>"100110",
1296=>"001111",
1312=>"011110",
1283=>"111100",
1286=>"111011",
1292=>"110101",
1304=>"101001",
1328=>"010001",
1315=>"100010",
1285=>"000111",
1290=>"001110",
1300=>"011100",
1320=>"111000",
1299=>"110011",
1318=>"100101",
1295=>"001001",
1310=>"010010",
1340=>"100100",
1339=>"001011",
1333=>"010110",
1321=>"101100",
1297=>"011011",
1314=>"110110",
1287=>"101111",
1294=>"011101",
1308=>"111010",
1336=>"110111",
1331=>"101101",
1317=>"011001",
1289=>"110010",
1298=>"100111",
1316=>"001101",
1291=>"011010",
1302=>"110100",
1324=>"101011",
1307=>"010101",
1334=>"101010",
1327=>"010111",
1309=>"101110",
1338=>"011111",
1335=>"111110",
1325=>"111111",
1305=>"111101",
1330=>"111001",
1319=>"110001",
1293=>"100001",
1306=>"000001",
1332=>"000010",
1323=>"000100",
1301=>"001000",
1322=>"010000",
1303=>"100000",
1326=>"000011",
1311=>"000110",
1342=>"001100",
1343=>"011000",
1341=>"110000",
1337=>"100011",
1329=>"000101",
1313=>"001010",
      
2561=>"101000",
2562=>"010011",
2564=>"100110",
2568=>"001111",
2576=>"011110",
2592=>"111100",
2563=>"111011",
2566=>"110101",
2572=>"101001",
2584=>"010001",
2608=>"100010",
2595=>"000111",
2565=>"001110",
2570=>"011100",
2580=>"111000",
2600=>"110011",
2579=>"100101",
2598=>"001001",
2575=>"010010",
2590=>"100100",
2620=>"001011",
2619=>"010110",
2613=>"101100",
2601=>"011011",
2577=>"110110",
2594=>"101111",
2567=>"011101",
2574=>"111010",
2588=>"110111",
2616=>"101101",
2611=>"011001",
2597=>"110010",
2569=>"100111",
2578=>"001101",
2596=>"011010",
2571=>"110100",
2582=>"101011",
2604=>"010101",
2587=>"101010",
2614=>"010111",
2607=>"101110",
2589=>"011111",
2618=>"111110",
2615=>"111111",
2605=>"111101",
2585=>"111001",
2610=>"110001",
2599=>"100001",
2573=>"000001",
2586=>"000010",
2612=>"000100",
2603=>"001000",
2581=>"010000",
2602=>"100000",
2583=>"000011",
2606=>"000110",
2591=>"001100",
2622=>"011000",
2623=>"110000",
2621=>"100011",
2617=>"000101",
2609=>"001010",
2593=>"010100",
      
1217=>"010011",
1218=>"100110",
1220=>"001111",
1224=>"011110",
1232=>"111100",
1248=>"111011",
1219=>"110101",
1222=>"101001",
1228=>"010001",
1240=>"100010",
1264=>"000111",
1251=>"001110",
1221=>"011100",
1226=>"111000",
1236=>"110011",
1256=>"100101",
1235=>"001001",
1254=>"010010",
1231=>"100100",
1246=>"001011",
1276=>"010110",
1275=>"101100",
1269=>"011011",
1257=>"110110",
1233=>"101111",
1250=>"011101",
1223=>"111010",
1230=>"110111",
1244=>"101101",
1272=>"011001",
1267=>"110010",
1253=>"100111",
1225=>"001101",
1234=>"011010",
1252=>"110100",
1227=>"101011",
1238=>"010101",
1260=>"101010",
1243=>"010111",
1270=>"101110",
1263=>"011111",
1245=>"111110",
1274=>"111111",
1271=>"111101",
1261=>"111001",
1241=>"110001",
1266=>"100001",
1255=>"000001",
1229=>"000010",
1242=>"000100",
1268=>"001000",
1259=>"010000",
1237=>"100000",
1258=>"000011",
1239=>"000110",
1262=>"001100",
1247=>"011000",
1278=>"110000",
1279=>"100011",
1277=>"000101",
1273=>"001010",
1265=>"010100",
1249=>"101000",
      
2433=>"100110",
2434=>"001111",
2436=>"011110",
2440=>"111100",
2448=>"111011",
2464=>"110101",
2435=>"101001",
2438=>"010001",
2444=>"100010",
2456=>"000111",
2480=>"001110",
2467=>"011100",
2437=>"111000",
2442=>"110011",
2452=>"100101",
2472=>"001001",
2451=>"010010",
2470=>"100100",
2447=>"001011",
2462=>"010110",
2492=>"101100",
2491=>"011011",
2485=>"110110",
2473=>"101111",
2449=>"011101",
2466=>"111010",
2439=>"110111",
2446=>"101101",
2460=>"011001",
2488=>"110010",
2483=>"100111",
2469=>"001101",
2441=>"011010",
2450=>"110100",
2468=>"101011",
2443=>"010101",
2454=>"101010",
2476=>"010111",
2459=>"101110",
2486=>"011111",
2479=>"111110",
2461=>"111111",
2490=>"111101",
2487=>"111001",
2477=>"110001",
2457=>"100001",
2482=>"000001",
2471=>"000010",
2445=>"000100",
2458=>"001000",
2484=>"010000",
2475=>"100000",
2453=>"000011",
2474=>"000110",
2455=>"001100",
2478=>"011000",
2463=>"110000",
2494=>"100011",
2495=>"000101",
2493=>"001010",
2489=>"010100",
2481=>"101000",
2465=>"010011",
      
961 =>"001111",
962 =>"011110",
964 =>"111100",
968 =>"111011",
976 =>"110101",
992 =>"101001",
963 =>"010001",
966 =>"100010",
972 =>"000111",
984 =>"001110",
1008=>"011100",
995 =>"111000",
965 =>"110011",
970 =>"100101",
980 =>"001001",
1000=>"010010",
979 =>"100100",
998 =>"001011",
975 =>"010110",
990 =>"101100",
1020=>"011011",
1019=>"110110",
1013=>"101111",
1001=>"011101",
977 =>"111010",
994 =>"110111",
967 =>"101101",
974 =>"011001",
988 =>"110010",
1016=>"100111",
1011=>"001101",
997 =>"011010",
969 =>"110100",
978 =>"101011",
996 =>"010101",
971 =>"101010",
982 =>"010111",
1004=>"101110",
987 =>"011111",
1014=>"111110",
1007=>"111111",
989 =>"111101",
1018=>"111001",
1015=>"110001",
1005=>"100001",
985 =>"000001",
1010=>"000010",
999 =>"000100",
973 =>"001000",
986 =>"010000",
1012=>"100000",
1003=>"000011",
981 =>"000110",
1002=>"001100",
983 =>"011000",
1006=>"110000",
991 =>"100011",
1022=>"000101",
1023=>"001010",
1021=>"010100",
1017=>"101000",
1009=>"010011",
993 =>"100110",
      
1921=>"011110",
1922=>"111100",
1924=>"111011",
1928=>"110101",
1936=>"101001",
1952=>"010001",
1923=>"100010",
1926=>"000111",
1932=>"001110",
1944=>"011100",
1968=>"111000",
1955=>"110011",
1925=>"100101",
1930=>"001001",
1940=>"010010",
1960=>"100100",
1939=>"001011",
1958=>"010110",
1935=>"101100",
1950=>"011011",
1980=>"110110",
1979=>"101111",
1973=>"011101",
1961=>"111010",
1937=>"110111",
1954=>"101101",
1927=>"011001",
1934=>"110010",
1948=>"100111",
1976=>"001101",
1971=>"011010",
1957=>"110100",
1929=>"101011",
1938=>"010101",
1956=>"101010",
1931=>"010111",
1942=>"101110",
1964=>"011111",
1947=>"111110",
1974=>"111111",
1967=>"111101",
1949=>"111001",
1978=>"110001",
1975=>"100001",
1965=>"000001",
1945=>"000010",
1970=>"000100",
1959=>"001000",
1933=>"010000",
1946=>"100000",
1972=>"000011",
1963=>"000110",
1941=>"001100",
1962=>"011000",
1943=>"110000",
1966=>"100011",
1951=>"000101",
1982=>"001010",
1983=>"010100",
1981=>"101000",
1977=>"010011",
1969=>"100110",
1953=>"001111",
      
3841=>"111100",
3842=>"111011",
3844=>"110101",
3848=>"101001",
3856=>"010001",
3872=>"100010",
3843=>"000111",
3846=>"001110",
3852=>"011100",
3864=>"111000",
3888=>"110011",
3875=>"100101",
3845=>"001001",
3850=>"010010",
3860=>"100100",
3880=>"001011",
3859=>"010110",
3878=>"101100",
3855=>"011011",
3870=>"110110",
3900=>"101111",
3899=>"011101",
3893=>"111010",
3881=>"110111",
3857=>"101101",
3874=>"011001",
3847=>"110010",
3854=>"100111",
3868=>"001101",
3896=>"011010",
3891=>"110100",
3877=>"101011",
3849=>"010101",
3858=>"101010",
3876=>"010111",
3851=>"101110",
3862=>"011111",
3884=>"111110",
3867=>"111111",
3894=>"111101",
3887=>"111001",
3869=>"110001",
3898=>"100001",
3895=>"000001",
3885=>"000010",
3865=>"000100",
3890=>"001000",
3879=>"010000",
3853=>"100000",
3866=>"000011",
3892=>"000110",
3883=>"001100",
3861=>"011000",
3882=>"110000",
3863=>"100011",
3886=>"000101",
3871=>"001010",
3902=>"010100",
3903=>"101000",
3901=>"010011",
3897=>"100110",
3889=>"001111",
3873=>"011110",
      
3777=>"111011",
3778=>"110101",
3780=>"101001",
3784=>"010001",
3792=>"100010",
3808=>"000111",
3779=>"001110",
3782=>"011100",
3788=>"111000",
3800=>"110011",
3824=>"100101",
3811=>"001001",
3781=>"010010",
3786=>"100100",
3796=>"001011",
3816=>"010110",
3795=>"101100",
3814=>"011011",
3791=>"110110",
3806=>"101111",
3836=>"011101",
3835=>"111010",
3829=>"110111",
3817=>"101101",
3793=>"011001",
3810=>"110010",
3783=>"100111",
3790=>"001101",
3804=>"011010",
3832=>"110100",
3827=>"101011",
3813=>"010101",
3785=>"101010",
3794=>"010111",
3812=>"101110",
3787=>"011111",
3798=>"111110",
3820=>"111111",
3803=>"111101",
3830=>"111001",
3823=>"110001",
3805=>"100001",
3834=>"000001",
3831=>"000010",
3821=>"000100",
3801=>"001000",
3826=>"010000",
3815=>"100000",
3789=>"000011",
3802=>"000110",
3828=>"001100",
3819=>"011000",
3797=>"110000",
3818=>"100011",
3799=>"000101",
3822=>"001010",
3807=>"010100",
3838=>"101000",
3839=>"010011",
3837=>"100110",
3833=>"001111",
3825=>"011110",
3809=>"111100",

3393=>"110101",
3394=>"101001",
3396=>"010001",
3400=>"100010",
3408=>"000111",
3424=>"001110",
3395=>"011100",
3398=>"111000",
3404=>"110011",
3416=>"100101",
3440=>"001001",
3427=>"010010",
3397=>"100100",
3402=>"001011",
3412=>"010110",
3432=>"101100",
3411=>"011011",
3430=>"110110",
3407=>"101111",
3422=>"011101",
3452=>"111010",
3451=>"110111",
3445=>"101101",
3433=>"011001",
3409=>"110010",
3426=>"100111",
3399=>"001101",
3406=>"011010",
3420=>"110100",
3448=>"101011",
3443=>"010101",
3429=>"101010",
3401=>"010111",
3410=>"101110",
3428=>"011111",
3403=>"111110",
3414=>"111111",
3436=>"111101",
3419=>"111001",
3446=>"110001",
3439=>"100001",
3421=>"000001",
3450=>"000010",
3447=>"000100",
3437=>"001000",
3417=>"010000",
3442=>"100000",
3431=>"000011",
3405=>"000110",
3418=>"001100",
3444=>"011000",
3435=>"110000",
3413=>"100011",
3434=>"000101",
3415=>"001010",
3438=>"010100",
3423=>"101000",
3454=>"010011",
3455=>"100110",
3453=>"001111",
3449=>"011110",
3441=>"111100",
3425=>"111011",

2625=>"101001",
2626=>"010001",
2628=>"100010",
2632=>"000111",
2640=>"001110",
2656=>"011100",
2627=>"111000",
2630=>"110011",
2636=>"100101",
2648=>"001001",
2672=>"010010",
2659=>"100100",
2629=>"001011",
2634=>"010110",
2644=>"101100",
2664=>"011011",
2643=>"110110",
2662=>"101111",
2639=>"011101",
2654=>"111010",
2684=>"110111",
2683=>"101101",
2677=>"011001",
2665=>"110010",
2641=>"100111",
2658=>"001101",
2631=>"011010",
2638=>"110100",
2652=>"101011",
2680=>"010101",
2675=>"101010",
2661=>"010111",
2633=>"101110",
2642=>"011111",
2660=>"111110",
2635=>"111111",
2646=>"111101",
2668=>"111001",
2651=>"110001",
2678=>"100001",
2671=>"000001",
2653=>"000010",
2682=>"000100",
2679=>"001000",
2669=>"010000",
2649=>"100000",
2674=>"000011",
2663=>"000110",
2637=>"001100",
2650=>"011000",
2676=>"110000",
2667=>"100011",
2645=>"000101",
2666=>"001010",
2647=>"010100",
2670=>"101000",
2655=>"010011",
2686=>"100110",
2687=>"001111",
2685=>"011110",
2681=>"111100",
2673=>"111011",
2657=>"110101",

1089=>"010001",
1090=>"100010",
1092=>"000111",
1096=>"001110",
1104=>"011100",
1120=>"111000",
1091=>"110011",
1094=>"100101",
1100=>"001001",
1112=>"010010",
1136=>"100100",
1123=>"001011",
1093=>"010110",
1098=>"101100",
1108=>"011011",
1128=>"110110",
1107=>"101111",
1126=>"011101",
1103=>"111010",
1118=>"110111",
1148=>"101101",
1147=>"011001",
1141=>"110010",
1129=>"100111",
1105=>"001101",
1122=>"011010",
1095=>"110100",
1102=>"101011",
1116=>"010101",
1144=>"101010",
1139=>"010111",
1125=>"101110",
1097=>"011111",
1106=>"111110",
1124=>"111111",
1099=>"111101",
1110=>"111001",
1132=>"110001",
1115=>"100001",
1142=>"000001",
1135=>"000010",
1117=>"000100",
1146=>"001000",
1143=>"010000",
1133=>"100000",
1113=>"000011",
1138=>"000110",
1127=>"001100",
1101=>"011000",
1114=>"110000",
1140=>"100011",
1131=>"000101",
1109=>"001010",
1130=>"010100",
1111=>"101000",
1134=>"010011",
1119=>"100110",
1150=>"001111",
1151=>"011110",
1149=>"111100",
1145=>"111011",
1137=>"110101",
1121=>"101001",

2177=>"100010",
2178=>"000111",
2180=>"001110",
2184=>"011100",
2192=>"111000",
2208=>"110011",
2179=>"100101",
2182=>"001001",
2188=>"010010",
2200=>"100100",
2224=>"001011",
2211=>"010110",
2181=>"101100",
2186=>"011011",
2196=>"110110",
2216=>"101111",
2195=>"011101",
2214=>"111010",
2191=>"110111",
2206=>"101101",
2236=>"011001",
2235=>"110010",
2229=>"100111",
2217=>"001101",
2193=>"011010",
2210=>"110100",
2183=>"101011",
2190=>"010101",
2204=>"101010",
2232=>"010111",
2227=>"101110",
2213=>"011111",
2185=>"111110",
2194=>"111111",
2212=>"111101",
2187=>"111001",
2198=>"110001",
2220=>"100001",
2203=>"000001",
2230=>"000010",
2223=>"000100",
2205=>"001000",
2234=>"010000",
2231=>"100000",
2221=>"000011",
2201=>"000110",
2226=>"001100",
2215=>"011000",
2189=>"110000",
2202=>"100011",
2228=>"000101",
2219=>"001010",
2197=>"010100",
2218=>"101000",
2199=>"010011",
2222=>"100110",
2207=>"001111",
2238=>"011110",
2239=>"111100",
2237=>"111011",
2233=>"110101",
2225=>"101001",
2209=>"010001",

449 =>"000111",
450 =>"001110",
452 =>"011100",
456 =>"111000",
464 =>"110011",
480 =>"100101",
451 =>"001001",
454 =>"010010",
460 =>"100100",
472 =>"001011",
496 =>"010110",
483 =>"101100",
453 =>"011011",
458 =>"110110",
468 =>"101111",
488 =>"011101",
467 =>"111010",
486 =>"110111",
463 =>"101101",
478 =>"011001",
508 =>"110010",
507 =>"100111",
501 =>"001101",
489 =>"011010",
465 =>"110100",
482 =>"101011",
455 =>"010101",
462 =>"101010",
476 =>"010111",
504 =>"101110",
499 =>"011111",
485 =>"111110",
457 =>"111111",
466 =>"111101",
484 =>"111001",
459 =>"110001",
470 =>"100001",
492 =>"000001",
475 =>"000010",
502 =>"000100",
495 =>"001000",
477 =>"010000",
506 =>"100000",
503 =>"000011",
493 =>"000110",
473 =>"001100",
498 =>"011000",
487 =>"110000",
461 =>"100011",
474 =>"000101",
500 =>"001010",
491 =>"010100",
469 =>"101000",
490 =>"010011",
471 =>"100110",
494 =>"001111",
479 =>"011110",
510 =>"111100",
511 =>"111011",
509 =>"110101",
505 =>"101001",
497 =>"010001",
481 =>"100010",

897 =>"001110",
898 =>"011100",
900 =>"111000",
904 =>"110011",
912 =>"100101",
928 =>"001001",
899 =>"010010",
902 =>"100100",
908 =>"001011",
920 =>"010110",
944 =>"101100",
931 =>"011011",
901 =>"110110",
906 =>"101111",
916 =>"011101",
936 =>"111010",
915 =>"110111",
934 =>"101101",
911 =>"011001",
926 =>"110010",
956 =>"100111",
955 =>"001101",
949 =>"011010",
937 =>"110100",
913 =>"101011",
930 =>"010101",
903 =>"101010",
910 =>"010111",
924 =>"101110",
952 =>"011111",
947 =>"111110",
933 =>"111111",
905 =>"111101",
914 =>"111001",
932 =>"110001",
907 =>"100001",
918 =>"000001",
940 =>"000010",
923 =>"000100",
950 =>"001000",
943 =>"010000",
925 =>"100000",
954 =>"000011",
951 =>"000110",
941 =>"001100",
921 =>"011000",
946 =>"110000",
935 =>"100011",
909 =>"000101",
922 =>"001010",
948 =>"010100",
939 =>"101000",
917 =>"010011",
938 =>"100110",
919 =>"001111",
942 =>"011110",
927 =>"111100",
958 =>"111011",
959 =>"110101",
957 =>"101001",
953 =>"010001",
945 =>"100010",
929 =>"000111",

1793=>"011100",
1794=>"111000",
1796=>"110011",
1800=>"100101",
1808=>"001001",
1824=>"010010",
1795=>"100100",
1798=>"001011",
1804=>"010110",
1816=>"101100",
1840=>"011011",
1827=>"110110",
1797=>"101111",
1802=>"011101",
1812=>"111010",
1832=>"110111",
1811=>"101101",
1830=>"011001",
1807=>"110010",
1822=>"100111",
1852=>"001101",
1851=>"011010",
1845=>"110100",
1833=>"101011",
1809=>"010101",
1826=>"101010",
1799=>"010111",
1806=>"101110",
1820=>"011111",
1848=>"111110",
1843=>"111111",
1829=>"111101",
1801=>"111001",
1810=>"110001",
1828=>"100001",
1803=>"000001",
1814=>"000010",
1836=>"000100",
1819=>"001000",
1846=>"010000",
1839=>"100000",
1821=>"000011",
1850=>"000110",
1847=>"001100",
1837=>"011000",
1817=>"110000",
1842=>"100011",
1831=>"000101",
1805=>"001010",
1818=>"010100",
1844=>"101000",
1835=>"010011",
1813=>"100110",
1834=>"001111",
1815=>"011110",
1838=>"111100",
1823=>"111011",
1854=>"110101",
1855=>"101001",
1853=>"010001",
1849=>"100010",
1841=>"000111",
1825=>"001110",
   
3585=>"111000",
3586=>"110011",
3588=>"100101",
3592=>"001001",
3600=>"010010",
3616=>"100100",
3587=>"001011",
3590=>"010110",
3596=>"101100",
3608=>"011011",
3632=>"110110",
3619=>"101111",
3589=>"011101",
3594=>"111010",
3604=>"110111",
3624=>"101101",
3603=>"011001",
3622=>"110010",
3599=>"100111",
3614=>"001101",
3644=>"011010",
3643=>"110100",
3637=>"101011",
3625=>"010101",
3601=>"101010",
3618=>"010111",
3591=>"101110",
3598=>"011111",
3612=>"111110",
3640=>"111111",
3635=>"111101",
3621=>"111001",
3593=>"110001",
3602=>"100001",
3620=>"000001",
3595=>"000010",
3606=>"000100",
3628=>"001000",
3611=>"010000",
3638=>"100000",
3631=>"000011",
3613=>"000110",
3642=>"001100",
3639=>"011000",
3629=>"110000",
3609=>"100011",
3634=>"000101",
3623=>"001010",
3597=>"010100",
3610=>"101000",
3636=>"010011",
3627=>"100110",
3605=>"001111",
3626=>"011110",
3607=>"111100",
3630=>"111011",
3615=>"110101",
3646=>"101001",
3647=>"010001",
3645=>"100010",
3641=>"000111",
3633=>"001110",
3617=>"011100",
   
3265=>"110011",
3266=>"100101",
3268=>"001001",
3272=>"010010",
3280=>"100100",
3296=>"001011",
3267=>"010110",
3270=>"101100",
3276=>"011011",
3288=>"110110",
3312=>"101111",
3299=>"011101",
3269=>"111010",
3274=>"110111",
3284=>"101101",
3304=>"011001",
3283=>"110010",
3302=>"100111",
3279=>"001101",
3294=>"011010",
3324=>"110100",
3323=>"101011",
3317=>"010101",
3305=>"101010",
3281=>"010111",
3298=>"101110",
3271=>"011111",
3278=>"111110",
3292=>"111111",
3320=>"111101",
3315=>"111001",
3301=>"110001",
3273=>"100001",
3282=>"000001",
3300=>"000010",
3275=>"000100",
3286=>"001000",
3308=>"010000",
3291=>"100000",
3318=>"000011",
3311=>"000110",
3293=>"001100",
3322=>"011000",
3319=>"110000",
3309=>"100011",
3289=>"000101",
3314=>"001010",
3303=>"010100",
3277=>"101000",
3290=>"010011",
3316=>"100110",
3307=>"001111",
3285=>"011110",
3306=>"111100",
3287=>"111011",
3310=>"110101",
3295=>"101001",
3326=>"010001",
3327=>"100010",
3325=>"000111",
3321=>"001110",
3313=>"011100",
3297=>"111000",
   
2369=>"100101",
2370=>"001001",
2372=>"010010",
2376=>"100100",
2384=>"001011",
2400=>"010110",
2371=>"101100",
2374=>"011011",
2380=>"110110",
2392=>"101111",
2416=>"011101",
2403=>"111010",
2373=>"110111",
2378=>"101101",
2388=>"011001",
2408=>"110010",
2387=>"100111",
2406=>"001101",
2383=>"011010",
2398=>"110100",
2428=>"101011",
2427=>"010101",
2421=>"101010",
2409=>"010111",
2385=>"101110",
2402=>"011111",
2375=>"111110",
2382=>"111111",
2396=>"111101",
2424=>"111001",
2419=>"110001",
2405=>"100001",
2377=>"000001",
2386=>"000010",
2404=>"000100",
2379=>"001000",
2390=>"010000",
2412=>"100000",
2395=>"000011",
2422=>"000110",
2415=>"001100",
2397=>"011000",
2426=>"110000",
2423=>"100011",
2413=>"000101",
2393=>"001010",
2418=>"010100",
2407=>"101000",
2381=>"010011",
2394=>"100110",
2420=>"001111",
2411=>"011110",
2389=>"111100",
2410=>"111011",
2391=>"110101",
2414=>"101001",
2399=>"010001",
2430=>"100010",
2431=>"000111",
2429=>"001110",
2425=>"011100",
2417=>"111000",
2401=>"110011",
   
577 =>"001001",
578 =>"010010",
580 =>"100100",
584 =>"001011",
592 =>"010110",
608 =>"101100",
579 =>"011011",
582 =>"110110",
588 =>"101111",
600 =>"011101",
624 =>"111010",
611 =>"110111",
581 =>"101101",
586 =>"011001",
596 =>"110010",
616 =>"100111",
595 =>"001101",
614 =>"011010",
591 =>"110100",
606 =>"101011",
636 =>"010101",
635 =>"101010",
629 =>"010111",
617 =>"101110",
593 =>"011111",
610 =>"111110",
583 =>"111111",
590 =>"111101",
604 =>"111001",
632 =>"110001",
627 =>"100001",
613 =>"000001",
585 =>"000010",
594 =>"000100",
612 =>"001000",
587 =>"010000",
598 =>"100000",
620 =>"000011",
603 =>"000110",
630 =>"001100",
623 =>"011000",
605 =>"110000",
634 =>"100011",
631 =>"000101",
621 =>"001010",
601 =>"010100",
626 =>"101000",
615 =>"010011",
589 =>"100110",
602 =>"001111",
628 =>"011110",
619 =>"111100",
597 =>"111011",
618 =>"110101",
599 =>"101001",
622 =>"010001",
607 =>"100010",
638 =>"000111",
639 =>"001110",
637 =>"011100",
633 =>"111000",
625 =>"110011",
609 =>"100101",
  
1153=>"010010",
1154=>"100100",
1156=>"001011",
1160=>"010110",
1168=>"101100",
1184=>"011011",
1155=>"110110",
1158=>"101111",
1164=>"011101",
1176=>"111010",
1200=>"110111",
1187=>"101101",
1157=>"011001",
1162=>"110010",
1172=>"100111",
1192=>"001101",
1171=>"011010",
1190=>"110100",
1167=>"101011",
1182=>"010101",
1212=>"101010",
1211=>"010111",
1205=>"101110",
1193=>"011111",
1169=>"111110",
1186=>"111111",
1159=>"111101",
1166=>"111001",
1180=>"110001",
1208=>"100001",
1203=>"000001",
1189=>"000010",
1161=>"000100",
1170=>"001000",
1188=>"010000",
1163=>"100000",
1174=>"000011",
1196=>"000110",
1179=>"001100",
1206=>"011000",
1199=>"110000",
1181=>"100011",
1210=>"000101",
1207=>"001010",
1197=>"010100",
1177=>"101000",
1202=>"010011",
1191=>"100110",
1165=>"001111",
1178=>"011110",
1204=>"111100",
1195=>"111011",
1173=>"110101",
1194=>"101001",
1175=>"010001",
1198=>"100010",
1183=>"000111",
1214=>"001110",
1215=>"011100",
1213=>"111000",
1209=>"110011",
1201=>"100101",
1185=>"001001",
    
2305=>"100100",
2306=>"001011",
2308=>"010110",
2312=>"101100",
2320=>"011011",
2336=>"110110",
2307=>"101111",
2310=>"011101",
2316=>"111010",
2328=>"110111",
2352=>"101101",
2339=>"011001",
2309=>"110010",
2314=>"100111",
2324=>"001101",
2344=>"011010",
2323=>"110100",
2342=>"101011",
2319=>"010101",
2334=>"101010",
2364=>"010111",
2363=>"101110",
2357=>"011111",
2345=>"111110",
2321=>"111111",
2338=>"111101",
2311=>"111001",
2318=>"110001",
2332=>"100001",
2360=>"000001",
2355=>"000010",
2341=>"000100",
2313=>"001000",
2322=>"010000",
2340=>"100000",
2315=>"000011",
2326=>"000110",
2348=>"001100",
2331=>"011000",
2358=>"110000",
2351=>"100011",
2333=>"000101",
2362=>"001010",
2359=>"010100",
2349=>"101000",
2329=>"010011",
2354=>"100110",
2343=>"001111",
2317=>"011110",
2330=>"111100",
2356=>"111011",
2347=>"110101",
2325=>"101001",
2346=>"010001",
2327=>"100010",
2350=>"000111",
2335=>"001110",
2366=>"011100",
2367=>"111000",
2365=>"110011",
2361=>"100101",
2353=>"001001",
2337=>"010010",
  
705 =>"001011",
706 =>"010110",
708 =>"101100",
712 =>"011011",
720 =>"110110",
736 =>"101111",
707 =>"011101",
710 =>"111010",
716 =>"110111",
728 =>"101101",
752 =>"011001",
739 =>"110010",
709 =>"100111",
714 =>"001101",
724 =>"011010",
744 =>"110100",
723 =>"101011",
742 =>"010101",
719 =>"101010",
734 =>"010111",
764 =>"101110",
763 =>"011111",
757 =>"111110",
745 =>"111111",
721 =>"111101",
738 =>"111001",
711 =>"110001",
718 =>"100001",
732 =>"000001",
760 =>"000010",
755 =>"000100",
741 =>"001000",
713 =>"010000",
722 =>"100000",
740 =>"000011",
715 =>"000110",
726 =>"001100",
748 =>"011000",
731 =>"110000",
758 =>"100011",
751 =>"000101",
733 =>"001010",
762 =>"010100",
759 =>"101000",
749 =>"010011",
729 =>"100110",
754 =>"001111",
743 =>"011110",
717 =>"111100",
730 =>"111011",
756 =>"110101",
747 =>"101001",
725 =>"010001",
746 =>"100010",
727 =>"000111",
750 =>"001110",
735 =>"011100",
766 =>"111000",
767 =>"110011",
765 =>"100101",
761 =>"001001",
753 =>"010010",
737 =>"100100",
  
1409=>"010110",
1410=>"101100",
1412=>"011011",
1416=>"110110",
1424=>"101111",
1440=>"011101",
1411=>"111010",
1414=>"110111",
1420=>"101101",
1432=>"011001",
1456=>"110010",
1443=>"100111",
1413=>"001101",
1418=>"011010",
1428=>"110100",
1448=>"101011",
1427=>"010101",
1446=>"101010",
1423=>"010111",
1438=>"101110",
1468=>"011111",
1467=>"111110",
1461=>"111111",
1449=>"111101",
1425=>"111001",
1442=>"110001",
1415=>"100001",
1422=>"000001",
1436=>"000010",
1464=>"000100",
1459=>"001000",
1445=>"010000",
1417=>"100000",
1426=>"000011",
1444=>"000110",
1419=>"001100",
1430=>"011000",
1452=>"110000",
1435=>"100011",
1462=>"000101",
1455=>"001010",
1437=>"010100",
1466=>"101000",
1463=>"010011",
1453=>"100110",
1433=>"001111",
1458=>"011110",
1447=>"111100",
1421=>"111011",
1434=>"110101",
1460=>"101001",
1451=>"010001",
1429=>"100010",
1450=>"000111",
1431=>"001110",
1454=>"011100",
1439=>"111000",
1470=>"110011",
1471=>"100101",
1469=>"001001",
1465=>"010010",
1457=>"100100",
1441=>"001011",
  
2817=>"101100",
2818=>"011011",
2820=>"110110",
2824=>"101111",
2832=>"011101",
2848=>"111010",
2819=>"110111",
2822=>"101101",
2828=>"011001",
2840=>"110010",
2864=>"100111",
2851=>"001101",
2821=>"011010",
2826=>"110100",
2836=>"101011",
2856=>"010101",
2835=>"101010",
2854=>"010111",
2831=>"101110",
2846=>"011111",
2876=>"111110",
2875=>"111111",
2869=>"111101",
2857=>"111001",
2833=>"110001",
2850=>"100001",
2823=>"000001",
2830=>"000010",
2844=>"000100",
2872=>"001000",
2867=>"010000",
2853=>"100000",
2825=>"000011",
2834=>"000110",
2852=>"001100",
2827=>"011000",
2838=>"110000",
2860=>"100011",
2843=>"000101",
2870=>"001010",
2863=>"010100",
2845=>"101000",
2874=>"010011",
2871=>"100110",
2861=>"001111",
2841=>"011110",
2866=>"111100",
2855=>"111011",
2829=>"110101",
2842=>"101001",
2868=>"010001",
2859=>"100010",
2837=>"000111",
2858=>"001110",
2839=>"011100",
2862=>"111000",
2847=>"110011",
2878=>"100101",
2879=>"001001",
2877=>"010010",
2873=>"100100",
2865=>"001011",
2849=>"010110",
  
1729=>"011011",
1730=>"110110",
1732=>"101111",
1736=>"011101",
1744=>"111010",
1760=>"110111",
1731=>"101101",
1734=>"011001",
1740=>"110010",
1752=>"100111",
1776=>"001101",
1763=>"011010",
1733=>"110100",
1738=>"101011",
1748=>"010101",
1768=>"101010",
1747=>"010111",
1766=>"101110",
1743=>"011111",
1758=>"111110",
1788=>"111111",
1787=>"111101",
1781=>"111001",
1769=>"110001",
1745=>"100001",
1762=>"000001",
1735=>"000010",
1742=>"000100",
1756=>"001000",
1784=>"010000",
1779=>"100000",
1765=>"000011",
1737=>"000110",
1746=>"001100",
1764=>"011000",
1739=>"110000",
1750=>"100011",
1772=>"000101",
1755=>"001010",
1782=>"010100",
1775=>"101000",
1757=>"010011",
1786=>"100110",
1783=>"001111",
1773=>"011110",
1753=>"111100",
1778=>"111011",
1767=>"110101",
1741=>"101001",
1754=>"010001",
1780=>"100010",
1771=>"000111",
1749=>"001110",
1770=>"011100",
1751=>"111000",
1774=>"110011",
1759=>"100101",
1790=>"001001",
1791=>"010010",
1789=>"100100",
1785=>"001011",
1777=>"010110",
1761=>"101100",
  
3457=>"110110",
3458=>"101111",
3460=>"011101",
3464=>"111010",
3472=>"110111",
3488=>"101101",
3459=>"011001",
3462=>"110010",
3468=>"100111",
3480=>"001101",
3504=>"011010",
3491=>"110100",
3461=>"101011",
3466=>"010101",
3476=>"101010",
3496=>"010111",
3475=>"101110",
3494=>"011111",
3471=>"111110",
3486=>"111111",
3516=>"111101",
3515=>"111001",
3509=>"110001",
3497=>"100001",
3473=>"000001",
3490=>"000010",
3463=>"000100",
3470=>"001000",
3484=>"010000",
3512=>"100000",
3507=>"000011",
3493=>"000110",
3465=>"001100",
3474=>"011000",
3492=>"110000",
3467=>"100011",
3478=>"000101",
3500=>"001010",
3483=>"010100",
3510=>"101000",
3503=>"010011",
3485=>"100110",
3514=>"001111",
3511=>"011110",
3501=>"111100",
3481=>"111011",
3506=>"110101",
3495=>"101001",
3469=>"010001",
3482=>"100010",
3508=>"000111",
3499=>"001110",
3477=>"011100",
3498=>"111000",
3479=>"110011",
3502=>"100101",
3487=>"001001",
3518=>"010010",
3519=>"100100",
3517=>"001011",
3513=>"010110",
3505=>"101100",
3489=>"011011",
  
3009=>"101111",
3010=>"011101",
3012=>"111010",
3016=>"110111",
3024=>"101101",
3040=>"011001",
3011=>"110010",
3014=>"100111",
3020=>"001101",
3032=>"011010",
3056=>"110100",
3043=>"101011",
3013=>"010101",
3018=>"101010",
3028=>"010111",
3048=>"101110",
3027=>"011111",
3046=>"111110",
3023=>"111111",
3038=>"111101",
3068=>"111001",
3067=>"110001",
3061=>"100001",
3049=>"000001",
3025=>"000010",
3042=>"000100",
3015=>"001000",
3022=>"010000",
3036=>"100000",
3064=>"000011",
3059=>"000110",
3045=>"001100",
3017=>"011000",
3026=>"110000",
3044=>"100011",
3019=>"000101",
3030=>"001010",
3052=>"010100",
3035=>"101000",
3062=>"010011",
3055=>"100110",
3037=>"001111",
3066=>"011110",
3063=>"111100",
3053=>"111011",
3033=>"110101",
3058=>"101001",
3047=>"010001",
3021=>"100010",
3034=>"000111",
3060=>"001110",
3051=>"011100",
3029=>"111000",
3050=>"110011",
3031=>"100101",
3054=>"001001",
3039=>"010010",
3070=>"100100",
3071=>"001011",
3069=>"010110",
3065=>"101100",
3057=>"011011",
3041=>"110110",
  
1857=>"011101",
1858=>"111010",
1860=>"110111",
1864=>"101101",
1872=>"011001",
1888=>"110010",
1859=>"100111",
1862=>"001101",
1868=>"011010",
1880=>"110100",
1904=>"101011",
1891=>"010101",
1861=>"101010",
1866=>"010111",
1876=>"101110",
1896=>"011111",
1875=>"111110",
1894=>"111111",
1871=>"111101",
1886=>"111001",
1916=>"110001",
1915=>"100001",
1909=>"000001",
1897=>"000010",
1873=>"000100",
1890=>"001000",
1863=>"010000",
1870=>"100000",
1884=>"000011",
1912=>"000110",
1907=>"001100",
1893=>"011000",
1865=>"110000",
1874=>"100011",
1892=>"000101",
1867=>"001010",
1878=>"010100",
1900=>"101000",
1883=>"010011",
1910=>"100110",
1903=>"001111",
1885=>"011110",
1914=>"111100",
1911=>"111011",
1901=>"110101",
1881=>"101001",
1906=>"010001",
1895=>"100010",
1869=>"000111",
1882=>"001110",
1908=>"011100",
1899=>"111000",
1877=>"110011",
1898=>"100101",
1879=>"001001",
1902=>"010010",
1887=>"100100",
1918=>"001011",
1919=>"010110",
1917=>"101100",
1913=>"011011",
1905=>"110110",
1889=>"101111",
  
3713=>"111010",
3714=>"110111",
3716=>"101101",
3720=>"011001",
3728=>"110010",
3744=>"100111",
3715=>"001101",
3718=>"011010",
3724=>"110100",
3736=>"101011",
3760=>"010101",
3747=>"101010",
3717=>"010111",
3722=>"101110",
3732=>"011111",
3752=>"111110",
3731=>"111111",
3750=>"111101",
3727=>"111001",
3742=>"110001",
3772=>"100001",
3771=>"000001",
3765=>"000010",
3753=>"000100",
3729=>"001000",
3746=>"010000",
3719=>"100000",
3726=>"000011",
3740=>"000110",
3768=>"001100",
3763=>"011000",
3749=>"110000",
3721=>"100011",
3730=>"000101",
3748=>"001010",
3723=>"010100",
3734=>"101000",
3756=>"010011",
3739=>"100110",
3766=>"001111",
3759=>"011110",
3741=>"111100",
3770=>"111011",
3767=>"110101",
3757=>"101001",
3737=>"010001",
3762=>"100010",
3751=>"000111",
3725=>"001110",
3738=>"011100",
3764=>"111000",
3755=>"110011",
3733=>"100101",
3754=>"001001",
3735=>"010010",
3758=>"100100",
3743=>"001011",
3774=>"010110",
3775=>"101100",
3773=>"011011",
3769=>"110110",
3761=>"101111",
3745=>"011101",
  
3521=>"110111",
3522=>"101101",
3524=>"011001",
3528=>"110010",
3536=>"100111",
3552=>"001101",
3523=>"011010",
3526=>"110100",
3532=>"101011",
3544=>"010101",
3568=>"101010",
3555=>"010111",
3525=>"101110",
3530=>"011111",
3540=>"111110",
3560=>"111111",
3539=>"111101",
3558=>"111001",
3535=>"110001",
3550=>"100001",
3580=>"000001",
3579=>"000010",
3573=>"000100",
3561=>"001000",
3537=>"010000",
3554=>"100000",
3527=>"000011",
3534=>"000110",
3548=>"001100",
3576=>"011000",
3571=>"110000",
3557=>"100011",
3529=>"000101",
3538=>"001010",
3556=>"010100",
3531=>"101000",
3542=>"010011",
3564=>"100110",
3547=>"001111",
3574=>"011110",
3567=>"111100",
3549=>"111011",
3578=>"110101",
3575=>"101001",
3565=>"010001",
3545=>"100010",
3570=>"000111",
3559=>"001110",
3533=>"011100",
3546=>"111000",
3572=>"110011",
3563=>"100101",
3541=>"001001",
3562=>"010010",
3543=>"100100",
3566=>"001011",
3551=>"010110",
3582=>"101100",
3583=>"011011",
3581=>"110110",
3577=>"101111",
3569=>"011101",
3553=>"111010",
  
2881=>"101101",
2882=>"011001",
2884=>"110010",
2888=>"100111",
2896=>"001101",
2912=>"011010",
2883=>"110100",
2886=>"101011",
2892=>"010101",
2904=>"101010",
2928=>"010111",
2915=>"101110",
2885=>"011111",
2890=>"111110",
2900=>"111111",
2920=>"111101",
2899=>"111001",
2918=>"110001",
2895=>"100001",
2910=>"000001",
2940=>"000010",
2939=>"000100",
2933=>"001000",
2921=>"010000",
2897=>"100000",
2914=>"000011",
2887=>"000110",
2894=>"001100",
2908=>"011000",
2936=>"110000",
2931=>"100011",
2917=>"000101",
2889=>"001010",
2898=>"010100",
2916=>"101000",
2891=>"010011",
2902=>"100110",
2924=>"001111",
2907=>"011110",
2934=>"111100",
2927=>"111011",
2909=>"110101",
2938=>"101001",
2935=>"010001",
2925=>"100010",
2905=>"000111",
2930=>"001110",
2919=>"011100",
2893=>"111000",
2906=>"110011",
2932=>"100101",
2923=>"001001",
2901=>"010010",
2922=>"100100",
2903=>"001011",
2926=>"010110",
2911=>"101100",
2942=>"011011",
2943=>"110110",
2941=>"101111",
2937=>"011101",
2929=>"111010",
2913=>"110111",
  
1601=>"011001",
1602=>"110010",
1604=>"100111",
1608=>"001101",
1616=>"011010",
1632=>"110100",
1603=>"101011",
1606=>"010101",
1612=>"101010",
1624=>"010111",
1648=>"101110",
1635=>"011111",
1605=>"111110",
1610=>"111111",
1620=>"111101",
1640=>"111001",
1619=>"110001",
1638=>"100001",
1615=>"000001",
1630=>"000010",
1660=>"000100",
1659=>"001000",
1653=>"010000",
1641=>"100000",
1617=>"000011",
1634=>"000110",
1607=>"001100",
1614=>"011000",
1628=>"110000",
1656=>"100011",
1651=>"000101",
1637=>"001010",
1609=>"010100",
1618=>"101000",
1636=>"010011",
1611=>"100110",
1622=>"001111",
1644=>"011110",
1627=>"111100",
1654=>"111011",
1647=>"110101",
1629=>"101001",
1658=>"010001",
1655=>"100010",
1645=>"000111",
1625=>"001110",
1650=>"011100",
1639=>"111000",
1613=>"110011",
1626=>"100101",
1652=>"001001",
1643=>"010010",
1621=>"100100",
1642=>"001011",
1623=>"010110",
1646=>"101100",
1631=>"011011",
1662=>"110110",
1663=>"101111",
1661=>"011101",
1657=>"111010",
1649=>"110111",
1633=>"101101",
  
3201=>"110010",
3202=>"100111",
3204=>"001101",
3208=>"011010",
3216=>"110100",
3232=>"101011",
3203=>"010101",
3206=>"101010",
3212=>"010111",
3224=>"101110",
3248=>"011111",
3235=>"111110",
3205=>"111111",
3210=>"111101",
3220=>"111001",
3240=>"110001",
3219=>"100001",
3238=>"000001",
3215=>"000010",
3230=>"000100",
3260=>"001000",
3259=>"010000",
3253=>"100000",
3241=>"000011",
3217=>"000110",
3234=>"001100",
3207=>"011000",
3214=>"110000",
3228=>"100011",
3256=>"000101",
3251=>"001010",
3237=>"010100",
3209=>"101000",
3218=>"010011",
3236=>"100110",
3211=>"001111",
3222=>"011110",
3244=>"111100",
3227=>"111011",
3254=>"110101",
3247=>"101001",
3229=>"010001",
3258=>"100010",
3255=>"000111",
3245=>"001110",
3225=>"011100",
3250=>"111000",
3239=>"110011",
3213=>"100101",
3226=>"001001",
3252=>"010010",
3243=>"100100",
3221=>"001011",
3242=>"010110",
3223=>"101100",
3246=>"011011",
3231=>"110110",
3262=>"101111",
3263=>"011101",
3261=>"111010",
3257=>"110111",
3249=>"101101",
3233=>"011001",
  
2497=>"100111",
2498=>"001101",
2500=>"011010",
2504=>"110100",
2512=>"101011",
2528=>"010101",
2499=>"101010",
2502=>"010111",
2508=>"101110",
2520=>"011111",
2544=>"111110",
2531=>"111111",
2501=>"111101",
2506=>"111001",
2516=>"110001",
2536=>"100001",
2515=>"000001",
2534=>"000010",
2511=>"000100",
2526=>"001000",
2556=>"010000",
2555=>"100000",
2549=>"000011",
2537=>"000110",
2513=>"001100",
2530=>"011000",
2503=>"110000",
2510=>"100011",
2524=>"000101",
2552=>"001010",
2547=>"010100",
2533=>"101000",
2505=>"010011",
2514=>"100110",
2532=>"001111",
2507=>"011110",
2518=>"111100",
2540=>"111011",
2523=>"110101",
2550=>"101001",
2543=>"010001",
2525=>"100010",
2554=>"000111",
2551=>"001110",
2541=>"011100",
2521=>"111000",
2546=>"110011",
2535=>"100101",
2509=>"001001",
2522=>"010010",
2548=>"100100",
2539=>"001011",
2517=>"010110",
2538=>"101100",
2519=>"011011",
2542=>"110110",
2527=>"101111",
2558=>"011101",
2559=>"111010",
2557=>"110111",
2553=>"101101",
2545=>"011001",
2529=>"110010",
  
833 =>"001101",
834 =>"011010",
836 =>"110100",
840 =>"101011",
848 =>"010101",
864 =>"101010",
835 =>"010111",
838 =>"101110",
844 =>"011111",
856 =>"111110",
880 =>"111111",
867 =>"111101",
837 =>"111001",
842 =>"110001",
852 =>"100001",
872 =>"000001",
851 =>"000010",
870 =>"000100",
847 =>"001000",
862 =>"010000",
892 =>"100000",
891 =>"000011",
885 =>"000110",
873 =>"001100",
849 =>"011000",
866 =>"110000",
839 =>"100011",
846 =>"000101",
860 =>"001010",
888 =>"010100",
883 =>"101000",
869 =>"010011",
841 =>"100110",
850 =>"001111",
868 =>"011110",
843 =>"111100",
854 =>"111011",
876 =>"110101",
859 =>"101001",
886 =>"010001",
879 =>"100010",
861 =>"000111",
890 =>"001110",
887 =>"011100",
877 =>"111000",
857 =>"110011",
882 =>"100101",
871 =>"001001",
845 =>"010010",
858 =>"100100",
884 =>"001011",
875 =>"010110",
853 =>"101100",
874 =>"011011",
855 =>"110110",
878 =>"101111",
863 =>"011101",
894 =>"111010",
895 =>"110111",
893 =>"101101",
889 =>"011001",
881 =>"110010",
865 =>"100111",
  
1665=>"011010",
1666=>"110100",
1668=>"101011",
1672=>"010101",
1680=>"101010",
1696=>"010111",
1667=>"101110",
1670=>"011111",
1676=>"111110",
1688=>"111111",
1712=>"111101",
1699=>"111001",
1669=>"110001",
1674=>"100001",
1684=>"000001",
1704=>"000010",
1683=>"000100",
1702=>"001000",
1679=>"010000",
1694=>"100000",
1724=>"000011",
1723=>"000110",
1717=>"001100",
1705=>"011000",
1681=>"110000",
1698=>"100011",
1671=>"000101",
1678=>"001010",
1692=>"010100",
1720=>"101000",
1715=>"010011",
1701=>"100110",
1673=>"001111",
1682=>"011110",
1700=>"111100",
1675=>"111011",
1686=>"110101",
1708=>"101001",
1691=>"010001",
1718=>"100010",
1711=>"000111",
1693=>"001110",
1722=>"011100",
1719=>"111000",
1709=>"110011",
1689=>"100101",
1714=>"001001",
1703=>"010010",
1677=>"100100",
1690=>"001011",
1716=>"010110",
1707=>"101100",
1685=>"011011",
1706=>"110110",
1687=>"101111",
1710=>"011101",
1695=>"111010",
1726=>"110111",
1727=>"101101",
1725=>"011001",
1721=>"110010",
1713=>"100111",
1697=>"001101",
  
3329=>"110100",
3330=>"101011",
3332=>"010101",
3336=>"101010",
3344=>"010111",
3360=>"101110",
3331=>"011111",
3334=>"111110",
3340=>"111111",
3352=>"111101",
3376=>"111001",
3363=>"110001",
3333=>"100001",
3338=>"000001",
3348=>"000010",
3368=>"000100",
3347=>"001000",
3366=>"010000",
3343=>"100000",
3358=>"000011",
3388=>"000110",
3387=>"001100",
3381=>"011000",
3369=>"110000",
3345=>"100011",
3362=>"000101",
3335=>"001010",
3342=>"010100",
3356=>"101000",
3384=>"010011",
3379=>"100110",
3365=>"001111",
3337=>"011110",
3346=>"111100",
3364=>"111011",
3339=>"110101",
3350=>"101001",
3372=>"010001",
3355=>"100010",
3382=>"000111",
3375=>"001110",
3357=>"011100",
3386=>"111000",
3383=>"110011",
3373=>"100101",
3353=>"001001",
3378=>"010010",
3367=>"100100",
3341=>"001011",
3354=>"010110",
3380=>"101100",
3371=>"011011",
3349=>"110110",
3370=>"101111",
3351=>"011101",
3374=>"111010",
3359=>"110111",
3390=>"101101",
3391=>"011001",
3389=>"110010",
3385=>"100111",
3377=>"001101",
3361=>"011010",
  
2753=>"101011",
2754=>"010101",
2756=>"101010",
2760=>"010111",
2768=>"101110",
2784=>"011111",
2755=>"111110",
2758=>"111111",
2764=>"111101",
2776=>"111001",
2800=>"110001",
2787=>"100001",
2757=>"000001",
2762=>"000010",
2772=>"000100",
2792=>"001000",
2771=>"010000",
2790=>"100000",
2767=>"000011",
2782=>"000110",
2812=>"001100",
2811=>"011000",
2805=>"110000",
2793=>"100011",
2769=>"000101",
2786=>"001010",
2759=>"010100",
2766=>"101000",
2780=>"010011",
2808=>"100110",
2803=>"001111",
2789=>"011110",
2761=>"111100",
2770=>"111011",
2788=>"110101",
2763=>"101001",
2774=>"010001",
2796=>"100010",
2779=>"000111",
2806=>"001110",
2799=>"011100",
2781=>"111000",
2810=>"110011",
2807=>"100101",
2797=>"001001",
2777=>"010010",
2802=>"100100",
2791=>"001011",
2765=>"010110",
2778=>"101100",
2804=>"011011",
2795=>"110110",
2773=>"101111",
2794=>"011101",
2775=>"111010",
2798=>"110111",
2783=>"101101",
2814=>"011001",
2815=>"110010",
2813=>"100111",
2809=>"001101",
2801=>"011010",
2785=>"110100",
  
1345=>"010101",
1346=>"101010",
1348=>"010111",
1352=>"101110",
1360=>"011111",
1376=>"111110",
1347=>"111111",
1350=>"111101",
1356=>"111001",
1368=>"110001",
1392=>"100001",
1379=>"000001",
1349=>"000010",
1354=>"000100",
1364=>"001000",
1384=>"010000",
1363=>"100000",
1382=>"000011",
1359=>"000110",
1374=>"001100",
1404=>"011000",
1403=>"110000",
1397=>"100011",
1385=>"000101",
1361=>"001010",
1378=>"010100",
1351=>"101000",
1358=>"010011",
1372=>"100110",
1400=>"001111",
1395=>"011110",
1381=>"111100",
1353=>"111011",
1362=>"110101",
1380=>"101001",
1355=>"010001",
1366=>"100010",
1388=>"000111",
1371=>"001110",
1398=>"011100",
1391=>"111000",
1373=>"110011",
1402=>"100101",
1399=>"001001",
1389=>"010010",
1369=>"100100",
1394=>"001011",
1383=>"010110",
1357=>"101100",
1370=>"011011",
1396=>"110110",
1387=>"101111",
1365=>"011101",
1386=>"111010",
1367=>"110111",
1390=>"101101",
1375=>"011001",
1406=>"110010",
1407=>"100111",
1405=>"001101",
1401=>"011010",
1393=>"110100",
1377=>"101011",
  
2689=>"101010",
2690=>"010111",
2692=>"101110",
2696=>"011111",
2704=>"111110",
2720=>"111111",
2691=>"111101",
2694=>"111001",
2700=>"110001",
2712=>"100001",
2736=>"000001",
2723=>"000010",
2693=>"000100",
2698=>"001000",
2708=>"010000",
2728=>"100000",
2707=>"000011",
2726=>"000110",
2703=>"001100",
2718=>"011000",
2748=>"110000",
2747=>"100011",
2741=>"000101",
2729=>"001010",
2705=>"010100",
2722=>"101000",
2695=>"010011",
2702=>"100110",
2716=>"001111",
2744=>"011110",
2739=>"111100",
2725=>"111011",
2697=>"110101",
2706=>"101001",
2724=>"010001",
2699=>"100010",
2710=>"000111",
2732=>"001110",
2715=>"011100",
2742=>"111000",
2735=>"110011",
2717=>"100101",
2746=>"001001",
2743=>"010010",
2733=>"100100",
2713=>"001011",
2738=>"010110",
2727=>"101100",
2701=>"011011",
2714=>"110110",
2740=>"101111",
2731=>"011101",
2709=>"111010",
2730=>"110111",
2711=>"101101",
2734=>"011001",
2719=>"110010",
2750=>"100111",
2751=>"001101",
2749=>"011010",
2745=>"110100",
2737=>"101011",
2721=>"010101",
  
1473=>"010111",
1474=>"101110",
1476=>"011111",
1480=>"111110",
1488=>"111111",
1504=>"111101",
1475=>"111001",
1478=>"110001",
1484=>"100001",
1496=>"000001",
1520=>"000010",
1507=>"000100",
1477=>"001000",
1482=>"010000",
1492=>"100000",
1512=>"000011",
1491=>"000110",
1510=>"001100",
1487=>"011000",
1502=>"110000",
1532=>"100011",
1531=>"000101",
1525=>"001010",
1513=>"010100",
1489=>"101000",
1506=>"010011",
1479=>"100110",
1486=>"001111",
1500=>"011110",
1528=>"111100",
1523=>"111011",
1509=>"110101",
1481=>"101001",
1490=>"010001",
1508=>"100010",
1483=>"000111",
1494=>"001110",
1516=>"011100",
1499=>"111000",
1526=>"110011",
1519=>"100101",
1501=>"001001",
1530=>"010010",
1527=>"100100",
1517=>"001011",
1497=>"010110",
1522=>"101100",
1511=>"011011",
1485=>"110110",
1498=>"101111",
1524=>"011101",
1515=>"111010",
1493=>"110111",
1514=>"101101",
1495=>"011001",
1518=>"110010",
1503=>"100111",
1534=>"001101",
1535=>"011010",
1533=>"110100",
1529=>"101011",
1521=>"010101",
1505=>"101010",
  
2945=>"101110",
2946=>"011111",
2948=>"111110",
2952=>"111111",
2960=>"111101",
2976=>"111001",
2947=>"110001",
2950=>"100001",
2956=>"000001",
2968=>"000010",
2992=>"000100",
2979=>"001000",
2949=>"010000",
2954=>"100000",
2964=>"000011",
2984=>"000110",
2963=>"001100",
2982=>"011000",
2959=>"110000",
2974=>"100011",
3004=>"000101",
3003=>"001010",
2997=>"010100",
2985=>"101000",
2961=>"010011",
2978=>"100110",
2951=>"001111",
2958=>"011110",
2972=>"111100",
3000=>"111011",
2995=>"110101",
2981=>"101001",
2953=>"010001",
2962=>"100010",
2980=>"000111",
2955=>"001110",
2966=>"011100",
2988=>"111000",
2971=>"110011",
2998=>"100101",
2991=>"001001",
2973=>"010010",
3002=>"100100",
2999=>"001011",
2989=>"010110",
2969=>"101100",
2994=>"011011",
2983=>"110110",
2957=>"101111",
2970=>"011101",
2996=>"111010",
2987=>"110111",
2965=>"101101",
2986=>"011001",
2967=>"110010",
2990=>"100111",
2975=>"001101",
3006=>"011010",
3007=>"110100",
3005=>"101011",
3001=>"010101",
2993=>"101010",
2977=>"010111",
  
1985=>"011111",
1986=>"111110",
1988=>"111111",
1992=>"111101",
2000=>"111001",
2016=>"110001",
1987=>"100001",
1990=>"000001",
1996=>"000010",
2008=>"000100",
2032=>"001000",
2019=>"010000",
1989=>"100000",
1994=>"000011",
2004=>"000110",
2024=>"001100",
2003=>"011000",
2022=>"110000",
1999=>"100011",
2014=>"000101",
2044=>"001010",
2043=>"010100",
2037=>"101000",
2025=>"010011",
2001=>"100110",
2018=>"001111",
1991=>"011110",
1998=>"111100",
2012=>"111011",
2040=>"110101",
2035=>"101001",
2021=>"010001",
1993=>"100010",
2002=>"000111",
2020=>"001110",
1995=>"011100",
2006=>"111000",
2028=>"110011",
2011=>"100101",
2038=>"001001",
2031=>"010010",
2013=>"100100",
2042=>"001011",
2039=>"010110",
2029=>"101100",
2009=>"011011",
2034=>"110110",
2023=>"101111",
1997=>"011101",
2010=>"111010",
2036=>"110111",
2027=>"101101",
2005=>"011001",
2026=>"110010",
2007=>"100111",
2030=>"001101",
2015=>"011010",
2046=>"110100",
2047=>"101011",
2045=>"010101",
2041=>"101010",
2033=>"010111",
2017=>"101110",
  
3969=>"111110",
3970=>"111111",
3972=>"111101",
3976=>"111001",
3984=>"110001",
4000=>"100001",
3971=>"000001",
3974=>"000010",
3980=>"000100",
3992=>"001000",
4016=>"010000",
4003=>"100000",
3973=>"000011",
3978=>"000110",
3988=>"001100",
4008=>"011000",
3987=>"110000",
4006=>"100011",
3983=>"000101",
3998=>"001010",
4028=>"010100",
4027=>"101000",
4021=>"010011",
4009=>"100110",
3985=>"001111",
4002=>"011110",
3975=>"111100",
3982=>"111011",
3996=>"110101",
4024=>"101001",
4019=>"010001",
4005=>"100010",
3977=>"000111",
3986=>"001110",
4004=>"011100",
3979=>"111000",
3990=>"110011",
4012=>"100101",
3995=>"001001",
4022=>"010010",
4015=>"100100",
3997=>"001011",
4026=>"010110",
4023=>"101100",
4013=>"011011",
3993=>"110110",
4018=>"101111",
4007=>"011101",
3981=>"111010",
3994=>"110111",
4020=>"101101",
4011=>"011001",
3989=>"110010",
4010=>"100111",
3991=>"001101",
4014=>"011010",
3999=>"110100",
4030=>"101011",
4031=>"010101",
4029=>"101010",
4025=>"010111",
4017=>"101110",
4001=>"011111",
  
4033=>"111111",
4034=>"111101",
4036=>"111001",
4040=>"110001",
4048=>"100001",
4064=>"000001",
4035=>"000010",
4038=>"000100",
4044=>"001000",
4056=>"010000",
4080=>"100000",
4067=>"000011",
4037=>"000110",
4042=>"001100",
4052=>"011000",
4072=>"110000",
4051=>"100011",
4070=>"000101",
4047=>"001010",
4062=>"010100",
4092=>"101000",
4091=>"010011",
4085=>"100110",
4073=>"001111",
4049=>"011110",
4066=>"111100",
4039=>"111011",
4046=>"110101",
4060=>"101001",
4088=>"010001",
4083=>"100010",
4069=>"000111",
4041=>"001110",
4050=>"011100",
4068=>"111000",
4043=>"110011",
4054=>"100101",
4076=>"001001",
4059=>"010010",
4086=>"100100",
4079=>"001011",
4061=>"010110",
4090=>"101100",
4087=>"011011",
4077=>"110110",
4057=>"101111",
4082=>"011101",
4071=>"111010",
4045=>"110111",
4058=>"101101",
4084=>"011001",
4075=>"110010",
4053=>"100111",
4074=>"001101",
4055=>"011010",
4078=>"110100",
4063=>"101011",
4094=>"010101",
4095=>"101010",
4093=>"010111",
4089=>"101110",
4081=>"011111",
4065=>"111110",
  
3905=>"111101",
3906=>"111001",
3908=>"110001",
3912=>"100001",
3920=>"000001",
3936=>"000010",
3907=>"000100",
3910=>"001000",
3916=>"010000",
3928=>"100000",
3952=>"000011",
3939=>"000110",
3909=>"001100",
3914=>"011000",
3924=>"110000",
3944=>"100011",
3923=>"000101",
3942=>"001010",
3919=>"010100",
3934=>"101000",
3964=>"010011",
3963=>"100110",
3957=>"001111",
3945=>"011110",
3921=>"111100",
3938=>"111011",
3911=>"110101",
3918=>"101001",
3932=>"010001",
3960=>"100010",
3955=>"000111",
3941=>"001110",
3913=>"011100",
3922=>"111000",
3940=>"110011",
3915=>"100101",
3926=>"001001",
3948=>"010010",
3931=>"100100",
3958=>"001011",
3951=>"010110",
3933=>"101100",
3962=>"011011",
3959=>"110110",
3949=>"101111",
3929=>"011101",
3954=>"111010",
3943=>"110111",
3917=>"101101",
3930=>"011001",
3956=>"110010",
3947=>"100111",
3925=>"001101",
3946=>"011010",
3927=>"110100",
3950=>"101011",
3935=>"010101",
3966=>"101010",
3967=>"010111",
3965=>"101110",
3961=>"011111",
3953=>"111110",
3937=>"111111",
  
3649=>"111001",
3650=>"110001",
3652=>"100001",
3656=>"000001",
3664=>"000010",
3680=>"000100",
3651=>"001000",
3654=>"010000",
3660=>"100000",
3672=>"000011",
3696=>"000110",
3683=>"001100",
3653=>"011000",
3658=>"110000",
3668=>"100011",
3688=>"000101",
3667=>"001010",
3686=>"010100",
3663=>"101000",
3678=>"010011",
3708=>"100110",
3707=>"001111",
3701=>"011110",
3689=>"111100",
3665=>"111011",
3682=>"110101",
3655=>"101001",
3662=>"010001",
3676=>"100010",
3704=>"000111",
3699=>"001110",
3685=>"011100",
3657=>"111000",
3666=>"110011",
3684=>"100101",
3659=>"001001",
3670=>"010010",
3692=>"100100",
3675=>"001011",
3702=>"010110",
3695=>"101100",
3677=>"011011",
3706=>"110110",
3703=>"101111",
3693=>"011101",
3673=>"111010",
3698=>"110111",
3687=>"101101",
3661=>"011001",
3674=>"110010",
3700=>"100111",
3691=>"001101",
3669=>"011010",
3690=>"110100",
3671=>"101011",
3694=>"010101",
3679=>"101010",
3710=>"010111",
3711=>"101110",
3709=>"011111",
3705=>"111110",
3697=>"111111",
3681=>"111101",
  
3137=>"110001",
3138=>"100001",
3140=>"000001",
3144=>"000010",
3152=>"000100",
3168=>"001000",
3139=>"010000",
3142=>"100000",
3148=>"000011",
3160=>"000110",
3184=>"001100",
3171=>"011000",
3141=>"110000",
3146=>"100011",
3156=>"000101",
3176=>"001010",
3155=>"010100",
3174=>"101000",
3151=>"010011",
3166=>"100110",
3196=>"001111",
3195=>"011110",
3189=>"111100",
3177=>"111011",
3153=>"110101",
3170=>"101001",
3143=>"010001",
3150=>"100010",
3164=>"000111",
3192=>"001110",
3187=>"011100",
3173=>"111000",
3145=>"110011",
3154=>"100101",
3172=>"001001",
3147=>"010010",
3158=>"100100",
3180=>"001011",
3163=>"010110",
3190=>"101100",
3183=>"011011",
3165=>"110110",
3194=>"101111",
3191=>"011101",
3181=>"111010",
3161=>"110111",
3186=>"101101",
3175=>"011001",
3149=>"110010",
3162=>"100111",
3188=>"001101",
3179=>"011010",
3157=>"110100",
3178=>"101011",
3159=>"010101",
3182=>"101010",
3167=>"010111",
3198=>"101110",
3199=>"011111",
3197=>"111110",
3193=>"111111",
3185=>"111101",
3169=>"111001",
  
2113=>"100001",
2114=>"000001",
2116=>"000010",
2120=>"000100",
2128=>"001000",
2144=>"010000",
2115=>"100000",
2118=>"000011",
2124=>"000110",
2136=>"001100",
2160=>"011000",
2147=>"110000",
2117=>"100011",
2122=>"000101",
2132=>"001010",
2152=>"010100",
2131=>"101000",
2150=>"010011",
2127=>"100110",
2142=>"001111",
2172=>"011110",
2171=>"111100",
2165=>"111011",
2153=>"110101",
2129=>"101001",
2146=>"010001",
2119=>"100010",
2126=>"000111",
2140=>"001110",
2168=>"011100",
2163=>"111000",
2149=>"110011",
2121=>"100101",
2130=>"001001",
2148=>"010010",
2123=>"100100",
2134=>"001011",
2156=>"010110",
2139=>"101100",
2166=>"011011",
2159=>"110110",
2141=>"101111",
2170=>"011101",
2167=>"111010",
2157=>"110111",
2137=>"101101",
2162=>"011001",
2151=>"110010",
2125=>"100111",
2138=>"001101",
2164=>"011010",
2155=>"110100",
2133=>"101011",
2154=>"010101",
2135=>"101010",
2158=>"010111",
2143=>"101110",
2174=>"011111",
2175=>"111110",
2173=>"111111",
2169=>"111101",
2161=>"111001",
2145=>"110001",

others=>"000000");
begin

process(clk)  begin
	if rising_edge(clk)  then
		if Rd = '1' then
			Data <= rom(conv_integer(addr));  -- First register
		end if;
	end if;
end process;
end Behavioral;

